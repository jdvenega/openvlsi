* NGSPICE file created from map9v3.ext - technology: scmos

* Black-box entry subcircuit for FILL abstract view
.subckt FILL gnd vdd
.ends

* Black-box entry subcircuit for BUFX2 abstract view
.subckt BUFX2 A gnd Y vdd
.ends

* Black-box entry subcircuit for NAND2X1 abstract view
.subckt NAND2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for INVX1 abstract view
.subckt INVX1 A gnd Y vdd
.ends

* Black-box entry subcircuit for DFFSR abstract view
.subckt DFFSR Q CLK R S D gnd vdd
.ends

* Black-box entry subcircuit for XOR2X1 abstract view
.subckt XOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for NOR2X1 abstract view
.subckt NOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for AOI21X1 abstract view
.subckt AOI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for NAND3X1 abstract view
.subckt NAND3X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for OAI21X1 abstract view
.subckt OAI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for NOR3X1 abstract view
.subckt NOR3X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for AND2X2 abstract view
.subckt AND2X2 A B gnd Y vdd
.ends

* Black-box entry subcircuit for AOI22X1 abstract view
.subckt AOI22X1 A B C D gnd Y vdd
.ends

* Black-box entry subcircuit for XNOR2X1 abstract view
.subckt XNOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for CLKBUF1 abstract view
.subckt CLKBUF1 A gnd Y vdd
.ends

* Black-box entry subcircuit for MUX2X1 abstract view
.subckt MUX2X1 A B S gnd Y vdd
.ends

.subckt map9v3 vdd gnd clock reset start N[0] N[1] N[2] N[3] N[4] N[5] N[6] N[7] N[8]
+ dp[0] dp[1] dp[2] dp[3] dp[4] dp[5] dp[6] dp[7] dp[8] done counter[0] counter[1]
+ counter[2] counter[3] counter[4] counter[5] counter[6] counter[7] sr[0] sr[1] sr[2]
+ sr[3] sr[4] sr[5] sr[6] sr[7]
XFILL_0_0_2 gnd vdd FILL
XFILL_1_1_0 gnd vdd FILL
XBUFX2_3 BUFX2_3/A gnd BUFX2_3/Y vdd BUFX2
XBUFX2_25 INVX1_15/A gnd dp[6] vdd BUFX2
XFILL_7_0_2 gnd vdd FILL
XNAND2X1_2 N[1] N[2] gnd INVX1_25/A vdd NAND2X1
XFILL_8_1_0 gnd vdd FILL
XINVX1_38 INVX1_38/A gnd DFFSR_3/D vdd INVX1
XDFFSR_19 BUFX2_31/A DFFSR_3/CLK BUFX2_9/Y vdd DFFSR_19/D gnd vdd DFFSR
XFILL_1_1_1 gnd vdd FILL
XBUFX2_26 BUFX2_26/A gnd dp[7] vdd BUFX2
XBUFX2_4 BUFX2_3/A gnd BUFX2_4/Y vdd BUFX2
XFILL_8_1_1 gnd vdd FILL
XNAND2X1_3 INVX1_26/Y NOR2X1_7/Y gnd INVX1_27/A vdd NAND2X1
XINVX1_39 reset gnd BUFX2_6/A vdd INVX1
XDFFSR_20 BUFX2_32/A CLKBUF1_1/Y BUFX2_9/Y vdd DFFSR_20/D gnd vdd DFFSR
XBUFX2_27 DFFSR_32/Q gnd dp[8] vdd BUFX2
XFILL_1_1_2 gnd vdd FILL
XXOR2X1_1 INVX1_27/A NOR2X1_1/B gnd XOR2X1_1/Y vdd XOR2X1
XNAND2X1_4 NAND2X1_4/A NAND2X1_4/B gnd DFFSR_9/D vdd NAND2X1
XBUFX2_5 BUFX2_6/A gnd BUFX2_5/Y vdd BUFX2
XFILL_8_1_2 gnd vdd FILL
XDFFSR_21 DFFSR_21/Q DFFSR_4/CLK DFFSR_4/R vdd DFFSR_21/D gnd vdd DFFSR
XBUFX2_6 BUFX2_6/A gnd DFFSR_4/R vdd BUFX2
XFILL_4_0_0 gnd vdd FILL
XBUFX2_28 DFFSR_16/Q gnd sr[0] vdd BUFX2
XNAND2X1_5 INVX1_25/A NOR2X1_10/Y gnd NAND3X1_4/B vdd NAND2X1
XDFFSR_22 BUFX2_34/A DFFSR_4/CLK DFFSR_4/R vdd DFFSR_22/D gnd vdd DFFSR
XFILL_4_0_1 gnd vdd FILL
XBUFX2_29 INVX1_8/A gnd sr[1] vdd BUFX2
XNAND2X1_6 INVX1_33/A NAND2X1_6/B gnd NAND2X1_6/Y vdd NAND2X1
XBUFX2_7 BUFX2_6/A gnd DFFSR_9/R vdd BUFX2
XDFFSR_23 DFFSR_23/Q DFFSR_4/CLK DFFSR_4/R vdd DFFSR_23/D gnd vdd DFFSR
XNOR2X1_1 BUFX2_13/A NOR2X1_1/B gnd NOR2X1_1/Y vdd NOR2X1
XFILL_4_0_2 gnd vdd FILL
XBUFX2_8 BUFX2_6/A gnd DFFSR_1/S vdd BUFX2
XBUFX2_30 BUFX2_30/A gnd sr[2] vdd BUFX2
XNAND2X1_7 NOR2X1_1/Y NOR2X1_2/Y gnd NOR2X1_14/B vdd NAND2X1
XFILL_5_1_0 gnd vdd FILL
XDFFSR_24 DFFSR_24/Q DFFSR_1/CLK DFFSR_1/S vdd DFFSR_24/D gnd vdd DFFSR
XNOR2X1_2 DFFSR_9/Q DFFSR_8/Q gnd NOR2X1_2/Y vdd NOR2X1
XBUFX2_9 BUFX2_6/A gnd BUFX2_9/Y vdd BUFX2
XBUFX2_31 BUFX2_31/A gnd sr[3] vdd BUFX2
XFILL_5_1_1 gnd vdd FILL
XDFFSR_25 INVX1_5/A DFFSR_3/CLK BUFX2_5/Y vdd DFFSR_25/D gnd vdd DFFSR
XBUFX2_32 BUFX2_32/A gnd sr[4] vdd BUFX2
XFILL_5_1_2 gnd vdd FILL
XNOR2X1_3 DFFSR_7/Q INVX1_4/Y gnd AND2X2_4/A vdd NOR2X1
XDFFSR_26 INVX1_7/A CLKBUF1_1/Y BUFX2_5/Y vdd MUX2X1_1/Y gnd vdd DFFSR
XFILL_1_0_0 gnd vdd FILL
XBUFX2_33 DFFSR_21/Q gnd sr[5] vdd BUFX2
XNOR2X1_4 DFFSR_16/Q MUX2X1_6/S gnd NOR2X1_4/Y vdd NOR2X1
XFILL_8_1 gnd vdd FILL
XDFFSR_27 INVX1_9/A DFFSR_3/CLK BUFX2_5/Y vdd MUX2X1_2/Y gnd vdd DFFSR
XFILL_8_0_0 gnd vdd FILL
XINVX1_10 BUFX2_30/A gnd INVX1_10/Y vdd INVX1
XFILL_1_0_1 gnd vdd FILL
XBUFX2_34 BUFX2_34/A gnd sr[6] vdd BUFX2
XAOI21X1_1 INVX1_5/Y MUX2X1_6/S NOR2X1_4/Y gnd DFFSR_25/D vdd AOI21X1
XNOR2X1_5 N[0] MUX2X1_6/S gnd NOR2X1_5/Y vdd NOR2X1
XFILL_8_0_1 gnd vdd FILL
XNAND3X1_1 NOR2X1_1/Y NOR2X1_2/Y NOR3X1_1/Y gnd OAI21X1_1/B vdd NAND3X1
XDFFSR_28 INVX1_11/A CLKBUF1_1/Y BUFX2_5/Y vdd MUX2X1_3/Y gnd vdd DFFSR
XINVX1_11 INVX1_11/A gnd MUX2X1_3/A vdd INVX1
XFILL_1_0_2 gnd vdd FILL
XFILL_2_1_0 gnd vdd FILL
XBUFX2_35 DFFSR_23/Q gnd sr[7] vdd BUFX2
XNOR2X1_6 NOR2X1_6/A NOR2X1_6/B gnd NOR2X1_6/Y vdd NOR2X1
XAOI21X1_2 INVX1_21/Y MUX2X1_6/S NOR2X1_5/Y gnd DFFSR_24/D vdd AOI21X1
XINVX1_12 BUFX2_31/A gnd INVX1_12/Y vdd INVX1
XFILL_9_1_0 gnd vdd FILL
XFILL_8_0_2 gnd vdd FILL
XDFFSR_29 INVX1_13/A CLKBUF1_1/Y BUFX2_5/Y vdd MUX2X1_4/Y gnd vdd DFFSR
XNAND3X1_2 DFFSR_3/Q INVX1_1/Y BUFX2_1/Y gnd MUX2X1_6/S vdd NAND3X1
XNOR2X1_7 DFFSR_8/Q BUFX2_3/Y gnd NOR2X1_7/Y vdd NOR2X1
XFILL_2_1_1 gnd vdd FILL
XAOI21X1_3 XNOR2X1_1/Y AOI21X1_3/B AOI21X1_3/C gnd NOR2X1_6/B vdd AOI21X1
XINVX1_1 INVX1_1/A gnd INVX1_1/Y vdd INVX1
XDFFSR_30 INVX1_15/A CLKBUF1_1/Y BUFX2_5/Y vdd MUX2X1_5/Y gnd vdd DFFSR
XNAND3X1_3 DFFSR_5/Q BUFX2_1/Y INVX1_23/Y gnd NAND3X1_3/Y vdd NAND3X1
XFILL_9_1_1 gnd vdd FILL
XINVX1_13 INVX1_13/A gnd INVX1_13/Y vdd INVX1
XNOR2X1_8 N[1] N[2] gnd NOR2X1_8/Y vdd NOR2X1
XOAI21X1_10 BUFX2_34/A BUFX2_4/Y INVX1_1/Y gnd AOI21X1_9/C vdd OAI21X1
XAOI21X1_4 BUFX2_2/Y INVX1_10/Y OAI21X1_5/Y gnd DFFSR_18/D vdd AOI21X1
XFILL_2_1_2 gnd vdd FILL
XINVX1_14 BUFX2_32/A gnd INVX1_14/Y vdd INVX1
XFILL_9_1_2 gnd vdd FILL
XINVX1_2 DFFSR_2/Q gnd INVX1_2/Y vdd INVX1
XDFFSR_31 BUFX2_26/A DFFSR_4/CLK DFFSR_4/R vdd DFFSR_31/D gnd vdd DFFSR
XNAND3X1_4 INVX1_1/A NAND3X1_4/B NAND3X1_4/C gnd NAND3X1_4/Y vdd NAND3X1
XNOR2X1_9 INVX1_26/Y NOR2X1_7/Y gnd NOR2X1_9/Y vdd NOR2X1
XFILL_3_1 gnd vdd FILL
XOAI21X1_11 DFFSR_16/Q BUFX2_2/Y INVX1_1/Y gnd AOI21X1_10/C vdd OAI21X1
XINVX1_3 DFFSR_5/Q gnd INVX1_3/Y vdd INVX1
XAOI21X1_5 BUFX2_1/Y INVX1_12/Y OAI21X1_6/Y gnd DFFSR_19/D vdd AOI21X1
XDFFSR_1 INVX1_1/A DFFSR_1/CLK vdd DFFSR_1/S DFFSR_1/D gnd vdd DFFSR
XDFFSR_32 DFFSR_32/Q DFFSR_4/CLK DFFSR_4/R vdd DFFSR_32/D gnd vdd DFFSR
XFILL_5_0_0 gnd vdd FILL
XINVX1_15 INVX1_15/A gnd INVX1_15/Y vdd INVX1
XNAND3X1_5 DFFSR_4/Q NOR2X1_1/Y NOR2X1_2/Y gnd AND2X2_2/B vdd NAND3X1
XOAI21X1_12 NOR2X1_7/Y AND2X2_1/Y INVX1_1/Y gnd OAI21X1_12/Y vdd OAI21X1
XFILL_3_2 gnd vdd FILL
XDFFSR_2 DFFSR_2/Q DFFSR_3/CLK BUFX2_9/Y vdd DFFSR_2/D gnd vdd DFFSR
XFILL_5_0_1 gnd vdd FILL
XAOI21X1_6 BUFX2_4/Y INVX1_14/Y OAI21X1_7/Y gnd DFFSR_20/D vdd AOI21X1
XINVX1_16 DFFSR_21/Q gnd INVX1_16/Y vdd INVX1
XINVX1_4 INVX1_4/A gnd INVX1_4/Y vdd INVX1
XNAND3X1_6 INVX1_25/A NOR2X1_10/Y NOR2X1_13/Y gnd INVX1_33/A vdd NAND3X1
XDFFSR_33 INVX1_22/A DFFSR_1/CLK DFFSR_1/S vdd DFFSR_33/D gnd vdd DFFSR
XOAI21X1_13 INVX1_1/Y INVX1_24/Y OAI21X1_12/Y gnd DFFSR_8/D vdd OAI21X1
XDFFSR_3 DFFSR_3/Q DFFSR_3/CLK BUFX2_9/Y vdd DFFSR_3/D gnd vdd DFFSR
XAOI21X1_7 BUFX2_1/Y INVX1_16/Y AOI21X1_7/C gnd DFFSR_21/D vdd AOI21X1
XINVX1_5 INVX1_5/A gnd INVX1_5/Y vdd INVX1
XINVX1_17 BUFX2_26/A gnd INVX1_17/Y vdd INVX1
XNOR3X1_1 NOR3X1_1/A NOR3X1_1/B BUFX2_16/A gnd NOR3X1_1/Y vdd NOR3X1
XFILL_5_0_2 gnd vdd FILL
XFILL_6_1_0 gnd vdd FILL
XNAND3X1_7 INVX1_31/Y INVX1_29/Y INVX1_35/Y gnd NOR2X1_14/A vdd NAND3X1
XAND2X2_1 BUFX2_3/Y DFFSR_8/Q gnd AND2X2_1/Y vdd AND2X2
XDFFSR_4 DFFSR_4/Q DFFSR_4/CLK DFFSR_4/R vdd DFFSR_4/D gnd vdd DFFSR
XOAI21X1_14 NOR2X1_8/Y INVX1_25/Y INVX1_1/A gnd NAND2X1_4/A vdd OAI21X1
XAOI21X1_8 BUFX2_3/Y MUX2X1_6/B AOI21X1_8/C gnd DFFSR_22/D vdd AOI21X1
XINVX1_6 DFFSR_4/Q gnd BUFX2_3/A vdd INVX1
XFILL_7_1 gnd vdd FILL
XINVX1_18 BUFX2_34/A gnd MUX2X1_6/B vdd INVX1
XNAND3X1_8 INVX1_31/Y INVX1_29/Y INVX1_30/Y gnd AOI22X1_2/D vdd NAND3X1
XFILL_6_1_1 gnd vdd FILL
XOAI21X1_15 NOR2X1_9/Y INVX1_27/Y INVX1_1/Y gnd NAND2X1_4/B vdd OAI21X1
XAND2X2_2 AND2X2_2/A AND2X2_2/B gnd AND2X2_2/Y vdd AND2X2
XAOI21X1_9 BUFX2_3/Y INVX1_20/Y AOI21X1_9/C gnd DFFSR_23/D vdd AOI21X1
XINVX1_7 INVX1_7/A gnd INVX1_7/Y vdd INVX1
XDFFSR_5 DFFSR_5/Q DFFSR_3/CLK BUFX2_9/Y vdd DFFSR_3/Q gnd vdd DFFSR
XINVX1_19 DFFSR_32/Q gnd MUX2X1_7/A vdd INVX1
XFILL_7_2 gnd vdd FILL
XFILL_6_1_2 gnd vdd FILL
XNAND3X1_9 INVX1_32/Y N[8] INVX1_33/Y gnd NAND3X1_9/Y vdd NAND3X1
XAND2X2_3 AND2X2_3/A AND2X2_3/B gnd DFFSR_15/D vdd AND2X2
XOAI21X1_16 N[3] INVX1_25/Y AOI21X1_12/Y gnd OAI21X1_17/C vdd OAI21X1
XFILL_7_3 gnd vdd FILL
XDFFSR_6 INVX1_4/A DFFSR_1/CLK DFFSR_1/S vdd start gnd vdd DFFSR
XINVX1_8 INVX1_8/A gnd INVX1_8/Y vdd INVX1
XFILL_2_0_0 gnd vdd FILL
XINVX1_20 DFFSR_23/Q gnd INVX1_20/Y vdd INVX1
XFILL_9_0_0 gnd vdd FILL
XOAI21X1_17 INVX1_1/A XOR2X1_1/Y OAI21X1_17/C gnd DFFSR_10/D vdd OAI21X1
XINVX1_9 INVX1_9/A gnd INVX1_9/Y vdd INVX1
XDFFSR_7 DFFSR_7/Q DFFSR_1/CLK DFFSR_1/S vdd INVX1_4/A gnd vdd DFFSR
XFILL_2_0_1 gnd vdd FILL
XAOI22X1_1 INVX1_1/A NAND2X1_6/Y AOI22X1_1/C AOI22X1_1/D gnd DFFSR_13/D vdd AOI22X1
XINVX1_21 DFFSR_24/Q gnd INVX1_21/Y vdd INVX1
XAND2X2_4 AND2X2_4/A DFFSR_2/Q gnd DFFSR_1/D vdd AND2X2
XXNOR2X1_1 DFFSR_21/Q DFFSR_23/Q gnd XNOR2X1_1/Y vdd XNOR2X1
XNOR2X1_10 N[3] N[4] gnd NOR2X1_10/Y vdd NOR2X1
XFILL_9_0_1 gnd vdd FILL
XDFFSR_8 DFFSR_8/Q DFFSR_9/CLK DFFSR_9/R vdd DFFSR_8/D gnd vdd DFFSR
XOAI21X1_18 N[3] INVX1_25/Y N[4] gnd NAND3X1_4/C vdd OAI21X1
XFILL_2_0_2 gnd vdd FILL
XFILL_3_1_0 gnd vdd FILL
XAOI22X1_2 DFFSR_4/Q NOR2X1_14/Y BUFX2_16/A AOI22X1_2/D gnd AOI22X1_2/Y vdd AOI22X1
XFILL_9_0_2 gnd vdd FILL
XINVX1_22 INVX1_22/A gnd INVX1_22/Y vdd INVX1
XXNOR2X1_2 BUFX2_31/A BUFX2_32/A gnd AOI21X1_3/B vdd XNOR2X1
XNOR2X1_11 INVX1_29/Y INVX1_30/Y gnd NOR2X1_11/Y vdd NOR2X1
XDFFSR_9 DFFSR_9/Q DFFSR_9/CLK DFFSR_9/R vdd DFFSR_9/D gnd vdd DFFSR
XBUFX2_10 DFFSR_8/Q gnd counter[0] vdd BUFX2
XOAI21X1_19 NOR2X1_1/B INVX1_27/A BUFX2_13/A gnd AND2X2_2/A vdd OAI21X1
XFILL_2_1 gnd vdd FILL
XINVX1_23 DFFSR_3/Q gnd INVX1_23/Y vdd INVX1
XFILL_3_1_1 gnd vdd FILL
XNOR2X1_12 NOR3X1_1/B AND2X2_2/B gnd NOR2X1_12/Y vdd NOR2X1
XBUFX2_11 DFFSR_9/Q gnd counter[1] vdd BUFX2
XOAI21X1_20 INVX1_1/A AND2X2_2/Y NAND3X1_4/Y gnd DFFSR_11/D vdd OAI21X1
XINVX1_24 N[1] gnd INVX1_24/Y vdd INVX1
XFILL_3_1_2 gnd vdd FILL
XNOR2X1_13 N[5] N[6] gnd NOR2X1_13/Y vdd NOR2X1
XBUFX2_12 NOR2X1_1/B gnd counter[2] vdd BUFX2
XOAI21X1_21 N[5] NAND3X1_4/B INVX1_1/A gnd OAI21X1_23/B vdd OAI21X1
XINVX1_25 INVX1_25/A gnd INVX1_25/Y vdd INVX1
XNOR2X1_14 NOR2X1_14/A NOR2X1_14/B gnd NOR2X1_14/Y vdd NOR2X1
XFILL_6_0_0 gnd vdd FILL
XBUFX2_13 BUFX2_13/A gnd counter[3] vdd BUFX2
XOAI21X1_22 NOR2X1_12/Y NOR2X1_11/Y INVX1_1/Y gnd OAI21X1_22/Y vdd OAI21X1
XAOI21X1_10 BUFX2_2/Y INVX1_8/Y AOI21X1_10/C gnd DFFSR_17/D vdd AOI21X1
XINVX1_26 DFFSR_9/Q gnd INVX1_26/Y vdd INVX1
XFILL_6_1 gnd vdd FILL
XCLKBUF1_1 clock gnd CLKBUF1_1/Y vdd CLKBUF1
XFILL_6_0_1 gnd vdd FILL
XBUFX2_14 NOR3X1_1/B gnd counter[4] vdd BUFX2
XAOI21X1_11 NAND3X1_3/Y INVX1_22/Y INVX1_1/A gnd DFFSR_33/D vdd AOI21X1
XINVX1_27 INVX1_27/A gnd INVX1_27/Y vdd INVX1
XCLKBUF1_2 clock gnd DFFSR_4/CLK vdd CLKBUF1
XOAI21X1_23 OAI21X1_23/A OAI21X1_23/B OAI21X1_22/Y gnd DFFSR_12/D vdd OAI21X1
XMUX2X1_1 INVX1_7/Y INVX1_8/Y MUX2X1_6/S gnd MUX2X1_1/Y vdd MUX2X1
XFILL_0_1_0 gnd vdd FILL
XFILL_6_2 gnd vdd FILL
XFILL_6_0_2 gnd vdd FILL
XFILL_7_1_0 gnd vdd FILL
XOAI21X1_1 BUFX2_17/A OAI21X1_1/B DFFSR_4/Q gnd NAND2X1_1/B vdd OAI21X1
XAOI21X1_12 INVX1_25/Y N[3] INVX1_1/Y gnd AOI21X1_12/Y vdd AOI21X1
XOAI21X1_24 N[5] NAND3X1_4/B N[6] gnd NAND2X1_6/B vdd OAI21X1
XBUFX2_15 NOR3X1_1/A gnd counter[5] vdd BUFX2
XCLKBUF1_3 clock gnd DFFSR_9/CLK vdd CLKBUF1
XINVX1_28 N[5] gnd INVX1_28/Y vdd INVX1
XMUX2X1_2 INVX1_9/Y INVX1_10/Y MUX2X1_6/S gnd MUX2X1_2/Y vdd MUX2X1
XFILL_0_1_1 gnd vdd FILL
XFILL_10_1 gnd vdd FILL
XFILL_7_1_1 gnd vdd FILL
XBUFX2_16 BUFX2_16/A gnd counter[6] vdd BUFX2
XAOI21X1_13 NOR2X1_10/Y INVX1_25/A INVX1_28/Y gnd OAI21X1_23/A vdd AOI21X1
XOAI21X1_2 INVX1_2/Y AND2X2_4/A INVX1_3/Y gnd DFFSR_2/D vdd OAI21X1
XOAI21X1_25 NOR3X1_1/B AND2X2_2/B NOR3X1_1/A gnd AOI22X1_1/C vdd OAI21X1
XCLKBUF1_4 clock gnd DFFSR_1/CLK vdd CLKBUF1
XMUX2X1_3 MUX2X1_3/A INVX1_12/Y MUX2X1_6/S gnd MUX2X1_3/Y vdd MUX2X1
XFILL_0_1_2 gnd vdd FILL
XDFFSR_10 NOR2X1_1/B DFFSR_9/CLK DFFSR_9/R vdd DFFSR_10/D gnd vdd DFFSR
XINVX1_29 NOR3X1_1/B gnd INVX1_29/Y vdd INVX1
XFILL_10_2 gnd vdd FILL
XFILL_7_1_2 gnd vdd FILL
XBUFX2_17 BUFX2_17/A gnd counter[7] vdd BUFX2
XOAI21X1_26 N[7] INVX1_33/A INVX1_1/A gnd INVX1_34/A vdd OAI21X1
XOAI21X1_3 XNOR2X1_1/Y AOI21X1_3/B DFFSR_4/Q gnd AOI21X1_3/C vdd OAI21X1
XAOI21X1_14 NOR2X1_12/Y INVX1_31/Y INVX1_1/A gnd AOI22X1_1/D vdd AOI21X1
XNAND3X1_10 INVX1_1/A OAI21X1_29/Y NAND3X1_9/Y gnd AND2X2_3/B vdd NAND3X1
XINVX1_30 AND2X2_2/B gnd INVX1_30/Y vdd INVX1
XMUX2X1_4 INVX1_13/Y INVX1_14/Y MUX2X1_6/S gnd MUX2X1_4/Y vdd MUX2X1
XCLKBUF1_5 clock gnd DFFSR_3/CLK vdd CLKBUF1
XDFFSR_11 BUFX2_13/A DFFSR_9/CLK DFFSR_9/R vdd DFFSR_11/D gnd vdd DFFSR
XFILL_3_0_0 gnd vdd FILL
XOAI21X1_4 DFFSR_4/Q DFFSR_16/Q INVX1_1/Y gnd NOR2X1_6/A vdd OAI21X1
XBUFX2_18 INVX1_22/A gnd done vdd BUFX2
XOAI21X1_27 INVX1_32/Y INVX1_33/Y INVX1_34/Y gnd OAI21X1_27/Y vdd OAI21X1
XMUX2X1_5 INVX1_15/Y INVX1_16/Y MUX2X1_6/S gnd MUX2X1_5/Y vdd MUX2X1
XFILL_1_1 gnd vdd FILL
XNAND3X1_11 DFFSR_4/Q INVX1_37/Y NOR2X1_14/Y gnd INVX1_38/A vdd NAND3X1
XINVX1_31 NOR3X1_1/A gnd INVX1_31/Y vdd INVX1
XDFFSR_12 NOR3X1_1/B DFFSR_1/CLK DFFSR_1/S vdd DFFSR_12/D gnd vdd DFFSR
XFILL_3_0_1 gnd vdd FILL
XOAI21X1_28 INVX1_1/A AOI22X1_2/Y OAI21X1_27/Y gnd DFFSR_14/D vdd OAI21X1
XBUFX2_19 DFFSR_24/Q gnd dp[0] vdd BUFX2
XOAI21X1_5 INVX1_8/A BUFX2_2/Y INVX1_1/Y gnd OAI21X1_5/Y vdd OAI21X1
XNAND3X1_12 INVX1_1/Y OAI21X1_30/Y INVX1_38/A gnd AND2X2_3/A vdd NAND3X1
XMUX2X1_6 INVX1_17/Y MUX2X1_6/B MUX2X1_6/S gnd DFFSR_31/D vdd MUX2X1
XINVX1_32 N[7] gnd INVX1_32/Y vdd INVX1
XFILL_3_0_2 gnd vdd FILL
XDFFSR_13 NOR3X1_1/A DFFSR_9/CLK DFFSR_9/R vdd DFFSR_13/D gnd vdd DFFSR
XFILL_4_1_0 gnd vdd FILL
XOAI21X1_6 BUFX2_30/A BUFX2_2/Y INVX1_1/Y gnd OAI21X1_6/Y vdd OAI21X1
XOAI21X1_29 N[7] INVX1_33/A INVX1_36/Y gnd OAI21X1_29/Y vdd OAI21X1
XMUX2X1_7 MUX2X1_7/A INVX1_20/Y MUX2X1_6/S gnd DFFSR_32/D vdd MUX2X1
XBUFX2_20 INVX1_5/A gnd dp[1] vdd BUFX2
XINVX1_33 INVX1_33/A gnd INVX1_33/Y vdd INVX1
XDFFSR_14 BUFX2_16/A DFFSR_9/CLK DFFSR_9/R vdd DFFSR_14/D gnd vdd DFFSR
XFILL_4_1_1 gnd vdd FILL
XOAI21X1_30 BUFX2_3/Y OAI21X1_1/B BUFX2_17/A gnd OAI21X1_30/Y vdd OAI21X1
XOAI21X1_7 BUFX2_31/A BUFX2_4/Y INVX1_1/Y gnd OAI21X1_7/Y vdd OAI21X1
XBUFX2_21 INVX1_7/A gnd dp[2] vdd BUFX2
XINVX1_34 INVX1_34/A gnd INVX1_34/Y vdd INVX1
XDFFSR_15 BUFX2_17/A DFFSR_9/CLK DFFSR_9/R vdd DFFSR_15/D gnd vdd DFFSR
XFILL_4_1_2 gnd vdd FILL
XOAI21X1_8 BUFX2_32/A BUFX2_1/Y INVX1_1/Y gnd AOI21X1_7/C vdd OAI21X1
XBUFX2_22 INVX1_9/A gnd dp[3] vdd BUFX2
XINVX1_35 BUFX2_16/A gnd INVX1_35/Y vdd INVX1
XDFFSR_16 DFFSR_16/Q DFFSR_4/CLK DFFSR_4/R vdd NOR2X1_6/Y gnd vdd DFFSR
XFILL_0_0_0 gnd vdd FILL
XOAI21X1_9 DFFSR_21/Q BUFX2_4/Y INVX1_1/Y gnd AOI21X1_8/C vdd OAI21X1
XBUFX2_23 INVX1_11/A gnd dp[4] vdd BUFX2
XFILL_7_0_0 gnd vdd FILL
XBUFX2_1 BUFX2_3/A gnd BUFX2_1/Y vdd BUFX2
XINVX1_36 N[8] gnd INVX1_36/Y vdd INVX1
XDFFSR_17 INVX1_8/A CLKBUF1_1/Y BUFX2_5/Y vdd DFFSR_17/D gnd vdd DFFSR
XFILL_0_0_1 gnd vdd FILL
XBUFX2_24 INVX1_13/A gnd dp[5] vdd BUFX2
XFILL_7_0_1 gnd vdd FILL
XBUFX2_2 BUFX2_3/A gnd BUFX2_2/Y vdd BUFX2
XINVX1_37 BUFX2_17/A gnd INVX1_37/Y vdd INVX1
XNAND2X1_1 INVX1_1/Y NAND2X1_1/B gnd DFFSR_4/D vdd NAND2X1
XDFFSR_18 BUFX2_30/A CLKBUF1_1/Y BUFX2_9/Y vdd DFFSR_18/D gnd vdd DFFSR
.ends

