magic
tech scmos
magscale 1 2
timestamp 1556508158
<< checkpaint >>
rect -76 -66 128 270
<< nwell >>
rect -16 96 68 210
<< ntransistor >>
rect 14 12 18 52
rect 30 12 34 52
rect 46 12 50 52
<< ptransistor >>
rect 14 108 18 188
rect 24 108 28 188
rect 40 148 44 188
<< ndiffusion >>
rect 4 51 14 52
rect 12 13 14 51
rect 4 12 14 13
rect 18 42 30 52
rect 18 14 20 42
rect 28 14 30 42
rect 18 12 30 14
rect 34 51 46 52
rect 34 13 36 51
rect 44 13 46 51
rect 34 12 46 13
rect 50 51 60 52
rect 50 13 52 51
rect 50 12 60 13
<< pdiffusion >>
rect 4 187 14 188
rect 12 109 14 187
rect 4 108 14 109
rect 18 108 24 188
rect 28 187 40 188
rect 28 109 30 187
rect 38 148 40 187
rect 44 187 54 188
rect 44 149 46 187
rect 44 148 54 149
rect 28 108 38 109
<< ndcontact >>
rect 4 13 12 51
rect 20 14 28 42
rect 36 13 44 51
rect 52 13 60 51
<< pdcontact >>
rect 4 109 12 187
rect 30 109 38 187
rect 46 149 54 187
<< psubstratepcontact >>
rect -4 -4 4 4
rect 28 -4 36 4
<< nsubstratencontact >>
rect -4 196 4 204
rect 28 196 36 204
<< polysilicon >>
rect 14 188 18 192
rect 24 188 28 192
rect 40 188 44 192
rect 40 130 44 148
rect 14 98 18 108
rect 24 106 28 108
rect 24 102 34 106
rect 8 94 18 98
rect 8 66 12 94
rect 30 86 34 102
rect 28 78 34 86
rect 14 52 18 62
rect 30 52 34 78
rect 46 52 50 126
rect 14 8 18 12
rect 30 8 34 12
rect 46 8 50 12
<< polycontact >>
rect 44 126 52 134
rect 20 78 28 86
rect 12 62 20 70
<< metal1 >>
rect -4 204 68 206
rect 4 196 28 204
rect 36 196 68 204
rect -4 194 68 196
rect 4 187 12 194
rect 4 108 12 109
rect 30 187 38 188
rect 46 187 54 194
rect 46 148 54 149
rect 46 114 52 126
rect 38 109 40 114
rect 30 108 40 109
rect 46 108 60 114
rect 20 86 28 94
rect 34 74 40 108
rect 52 106 60 108
rect 4 72 12 74
rect 4 70 20 72
rect 4 66 12 70
rect 34 66 60 74
rect 6 52 42 56
rect 52 52 58 66
rect 4 51 44 52
rect 12 50 36 51
rect 4 12 12 13
rect 20 42 28 44
rect 20 6 28 14
rect 36 12 44 13
rect 52 51 60 52
rect 52 12 60 13
rect -4 4 68 6
rect 4 -4 28 4
rect 36 -4 68 4
rect -4 -6 68 -4
<< m1p >>
rect 52 106 60 114
rect 20 86 28 94
rect 4 66 12 74
rect 52 66 60 74
<< labels >>
rlabel metal1 8 0 8 0 4 gnd
rlabel metal1 8 200 8 200 4 vdd
rlabel metal1 8 70 8 70 4 A
rlabel metal1 24 90 24 90 4 B
rlabel metal1 56 70 56 70 4 Y
rlabel metal1 56 110 56 110 4 C
<< properties >>
string path 26.000 33.000 30.000 33.000 30.000 37.000 26.000 37.000 26.000 33.000 
<< end >>
