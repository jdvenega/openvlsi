VERSION 5.3 ;
   NAMESCASESENSITIVE ON ;
   NOWIREEXTENSIONATPIN ON ;
   DIVIDERCHAR "/" ;
   BUSBITCHARS "[]" ;
UNITS
   DATABASE MICRONS 1000 ;
END UNITS

MACRO map9v3
   CLASS BLOCK ;
   FOREIGN map9v3 ;
   ORIGIN 1.9000 4.0000 ;
   SIZE 231.0000 BY 208.3000 ;
   PIN vdd
      PORT
         LAYER metal1 ;
	    RECT 0.4000 200.4000 226.8000 201.6000 ;
	    RECT 2.8000 193.0000 3.6000 200.4000 ;
	    RECT 6.0000 195.8000 6.8000 200.4000 ;
	    RECT 9.2000 195.8000 10.0000 200.4000 ;
	    RECT 12.4000 195.8000 13.2000 200.4000 ;
	    RECT 15.6000 195.8000 16.4000 200.4000 ;
	    RECT 23.6000 195.8000 24.4000 200.4000 ;
	    RECT 26.8000 195.8000 27.6000 200.4000 ;
	    RECT 33.2000 195.8000 34.0000 200.4000 ;
	    RECT 36.4000 195.8000 37.2000 200.4000 ;
	    RECT 39.6000 195.8000 40.4000 200.4000 ;
	    RECT 42.8000 193.0000 43.6000 200.4000 ;
	    RECT 50.8000 195.8000 51.6000 200.4000 ;
	    RECT 54.0000 195.8000 54.8000 200.4000 ;
	    RECT 57.2000 195.8000 58.0000 200.4000 ;
	    RECT 60.4000 195.8000 61.2000 200.4000 ;
	    RECT 68.4000 195.8000 69.2000 200.4000 ;
	    RECT 71.6000 195.8000 72.4000 200.4000 ;
	    RECT 78.0000 195.8000 78.8000 200.4000 ;
	    RECT 81.2000 195.8000 82.0000 200.4000 ;
	    RECT 84.4000 195.8000 85.2000 200.4000 ;
	    RECT 87.6000 193.0000 88.4000 200.4000 ;
	    RECT 92.4000 193.0000 93.2000 200.4000 ;
	    RECT 97.2000 193.0000 98.0000 200.4000 ;
	    RECT 100.4000 195.8000 101.2000 200.4000 ;
	    RECT 105.2000 193.0000 106.0000 200.4000 ;
	    RECT 33.0000 191.8000 33.8000 192.0000 ;
	    RECT 36.4000 191.8000 37.2000 192.4000 ;
	    RECT 77.8000 191.8000 78.6000 192.0000 ;
	    RECT 81.2000 191.8000 82.0000 192.4000 ;
	    RECT 113.2000 191.8000 114.0000 200.4000 ;
	    RECT 114.8000 195.8000 115.6000 200.4000 ;
	    RECT 118.0000 195.8000 118.8000 200.4000 ;
	    RECT 121.2000 195.8000 122.0000 200.4000 ;
	    RECT 127.6000 195.8000 128.4000 200.4000 ;
	    RECT 130.8000 195.8000 131.6000 200.4000 ;
	    RECT 138.8000 195.8000 139.6000 200.4000 ;
	    RECT 142.0000 195.8000 142.8000 200.4000 ;
	    RECT 145.2000 195.8000 146.0000 200.4000 ;
	    RECT 148.4000 195.8000 149.2000 200.4000 ;
	    RECT 150.0000 195.8000 150.8000 200.4000 ;
	    RECT 153.2000 196.2000 154.0000 200.4000 ;
	    RECT 162.8000 193.0000 163.6000 200.4000 ;
	    RECT 166.0000 195.8000 166.8000 200.4000 ;
	    RECT 169.2000 195.8000 170.0000 200.4000 ;
	    RECT 172.4000 195.8000 173.2000 200.4000 ;
	    RECT 175.6000 195.8000 176.4000 200.4000 ;
	    RECT 183.6000 195.8000 184.4000 200.4000 ;
	    RECT 186.8000 195.8000 187.6000 200.4000 ;
	    RECT 193.2000 195.8000 194.0000 200.4000 ;
	    RECT 196.4000 195.8000 197.2000 200.4000 ;
	    RECT 199.6000 195.8000 200.4000 200.4000 ;
	    RECT 118.0000 191.8000 118.8000 192.4000 ;
	    RECT 121.2000 191.8000 122.2000 192.0000 ;
	    RECT 193.0000 191.8000 193.8000 192.0000 ;
	    RECT 196.4000 191.8000 197.2000 192.4000 ;
	    RECT 201.2000 191.8000 202.0000 200.4000 ;
	    RECT 209.2000 193.0000 210.0000 200.4000 ;
	    RECT 214.0000 195.8000 214.8000 200.4000 ;
	    RECT 217.2000 193.0000 218.0000 200.4000 ;
	    RECT 222.0000 195.8000 222.8000 200.4000 ;
	    RECT 10.2000 191.2000 37.2000 191.8000 ;
	    RECT 55.0000 191.2000 82.0000 191.8000 ;
	    RECT 118.0000 191.2000 145.0000 191.8000 ;
	    RECT 10.2000 191.0000 11.0000 191.2000 ;
	    RECT 55.0000 191.0000 55.8000 191.2000 ;
	    RECT 144.2000 191.0000 145.0000 191.2000 ;
	    RECT 170.2000 191.2000 197.2000 191.8000 ;
	    RECT 170.2000 191.0000 171.0000 191.2000 ;
	    RECT 23.0000 170.8000 23.8000 171.0000 ;
	    RECT 91.8000 170.8000 92.6000 171.0000 ;
	    RECT 160.6000 170.8000 161.4000 171.0000 ;
	    RECT 221.0000 170.8000 221.8000 171.0000 ;
	    RECT 23.0000 170.2000 50.0000 170.8000 ;
	    RECT 91.8000 170.2000 118.8000 170.8000 ;
	    RECT 160.6000 170.2000 187.6000 170.8000 ;
	    RECT 2.8000 161.6000 3.6000 169.0000 ;
	    RECT 6.0000 161.6000 6.8000 166.2000 ;
	    RECT 10.4000 161.6000 11.2000 170.2000 ;
	    RECT 45.8000 170.0000 46.8000 170.2000 ;
	    RECT 15.6000 161.6000 16.4000 169.8000 ;
	    RECT 49.2000 169.6000 50.0000 170.2000 ;
	    RECT 18.8000 161.6000 19.6000 166.2000 ;
	    RECT 22.0000 161.6000 22.8000 166.2000 ;
	    RECT 25.2000 161.6000 26.0000 166.2000 ;
	    RECT 28.4000 161.6000 29.2000 166.2000 ;
	    RECT 36.4000 161.6000 37.2000 166.2000 ;
	    RECT 39.6000 161.6000 40.4000 166.2000 ;
	    RECT 46.0000 161.6000 46.8000 166.2000 ;
	    RECT 49.2000 161.6000 50.0000 166.2000 ;
	    RECT 52.4000 161.6000 53.2000 166.2000 ;
	    RECT 54.0000 161.6000 54.8000 166.2000 ;
	    RECT 57.2000 161.6000 58.0000 166.2000 ;
	    RECT 66.4000 161.6000 67.2000 170.2000 ;
	    RECT 71.6000 161.6000 72.4000 169.8000 ;
	    RECT 76.4000 161.6000 77.2000 169.0000 ;
	    RECT 81.2000 161.6000 82.0000 170.2000 ;
	    RECT 114.6000 170.0000 115.6000 170.2000 ;
	    RECT 118.0000 169.6000 118.8000 170.2000 ;
	    RECT 85.4000 161.6000 86.2000 166.2000 ;
	    RECT 87.6000 161.6000 88.4000 166.2000 ;
	    RECT 90.8000 161.6000 91.6000 166.2000 ;
	    RECT 94.0000 161.6000 94.8000 166.2000 ;
	    RECT 97.2000 161.6000 98.0000 166.2000 ;
	    RECT 105.2000 161.6000 106.0000 166.2000 ;
	    RECT 108.4000 161.6000 109.2000 166.2000 ;
	    RECT 114.8000 161.6000 115.6000 166.2000 ;
	    RECT 118.0000 161.6000 118.8000 166.2000 ;
	    RECT 121.2000 161.6000 122.0000 166.2000 ;
	    RECT 124.4000 161.6000 125.2000 169.0000 ;
	    RECT 129.2000 161.6000 130.0000 169.8000 ;
	    RECT 134.4000 161.6000 135.2000 170.2000 ;
	    RECT 138.8000 161.6000 139.6000 166.2000 ;
	    RECT 142.0000 161.6000 142.8000 166.2000 ;
	    RECT 143.6000 161.6000 144.4000 170.2000 ;
	    RECT 183.4000 170.0000 184.2000 170.2000 ;
	    RECT 186.8000 169.6000 187.6000 170.2000 ;
	    RECT 194.8000 170.2000 221.8000 170.8000 ;
	    RECT 194.8000 169.6000 195.6000 170.2000 ;
	    RECT 198.2000 170.0000 199.0000 170.2000 ;
	    RECT 150.0000 161.6000 150.8000 166.2000 ;
	    RECT 156.4000 161.6000 157.2000 166.2000 ;
	    RECT 159.6000 161.6000 160.4000 166.2000 ;
	    RECT 162.8000 161.6000 163.6000 166.2000 ;
	    RECT 166.0000 161.6000 166.8000 166.2000 ;
	    RECT 174.0000 161.6000 174.8000 166.2000 ;
	    RECT 177.2000 161.6000 178.0000 166.2000 ;
	    RECT 183.6000 161.6000 184.4000 166.2000 ;
	    RECT 186.8000 161.6000 187.6000 166.2000 ;
	    RECT 190.0000 161.6000 190.8000 166.2000 ;
	    RECT 191.6000 161.6000 192.4000 166.2000 ;
	    RECT 194.8000 161.6000 195.6000 166.2000 ;
	    RECT 198.0000 161.6000 198.8000 166.2000 ;
	    RECT 204.4000 161.6000 205.2000 166.2000 ;
	    RECT 207.6000 161.6000 208.4000 166.2000 ;
	    RECT 215.6000 161.6000 216.4000 166.2000 ;
	    RECT 218.8000 161.6000 219.6000 166.2000 ;
	    RECT 222.0000 161.6000 222.8000 166.2000 ;
	    RECT 225.2000 161.6000 226.0000 166.2000 ;
	    RECT 0.4000 160.4000 226.8000 161.6000 ;
	    RECT 2.8000 153.0000 3.6000 160.4000 ;
	    RECT 6.0000 155.8000 6.8000 160.4000 ;
	    RECT 9.2000 155.8000 10.0000 160.4000 ;
	    RECT 12.4000 155.8000 13.2000 160.4000 ;
	    RECT 15.6000 155.8000 16.4000 160.4000 ;
	    RECT 23.6000 155.8000 24.4000 160.4000 ;
	    RECT 26.8000 155.8000 27.6000 160.4000 ;
	    RECT 33.2000 155.8000 34.0000 160.4000 ;
	    RECT 36.4000 155.8000 37.2000 160.4000 ;
	    RECT 39.6000 155.8000 40.4000 160.4000 ;
	    RECT 41.8000 155.8000 42.6000 160.4000 ;
	    RECT 33.0000 151.8000 33.8000 152.0000 ;
	    RECT 36.4000 151.8000 37.2000 152.4000 ;
	    RECT 46.0000 151.8000 46.8000 160.4000 ;
	    RECT 50.8000 153.0000 51.6000 160.4000 ;
	    RECT 54.0000 155.8000 54.8000 160.4000 ;
	    RECT 62.0000 155.8000 62.8000 160.4000 ;
	    RECT 65.2000 155.8000 66.0000 160.4000 ;
	    RECT 68.4000 155.8000 69.2000 160.4000 ;
	    RECT 74.8000 155.8000 75.6000 160.4000 ;
	    RECT 78.0000 155.8000 78.8000 160.4000 ;
	    RECT 86.0000 155.8000 86.8000 160.4000 ;
	    RECT 89.2000 155.8000 90.0000 160.4000 ;
	    RECT 92.4000 155.8000 93.2000 160.4000 ;
	    RECT 95.6000 155.8000 96.4000 160.4000 ;
	    RECT 97.2000 155.8000 98.0000 160.4000 ;
	    RECT 100.4000 155.8000 101.2000 160.4000 ;
	    RECT 103.6000 155.8000 104.4000 160.4000 ;
	    RECT 110.0000 155.8000 110.8000 160.4000 ;
	    RECT 113.2000 155.8000 114.0000 160.4000 ;
	    RECT 121.2000 155.8000 122.0000 160.4000 ;
	    RECT 124.4000 155.8000 125.2000 160.4000 ;
	    RECT 127.6000 155.8000 128.4000 160.4000 ;
	    RECT 130.8000 155.8000 131.6000 160.4000 ;
	    RECT 133.0000 155.8000 133.8000 160.4000 ;
	    RECT 65.2000 151.8000 66.0000 152.4000 ;
	    RECT 68.6000 151.8000 69.4000 152.0000 ;
	    RECT 100.4000 151.8000 101.2000 152.4000 ;
	    RECT 103.6000 151.8000 104.6000 152.0000 ;
	    RECT 137.2000 151.8000 138.0000 160.4000 ;
	    RECT 140.4000 155.8000 141.2000 160.4000 ;
	    RECT 143.6000 155.8000 144.4000 160.4000 ;
	    RECT 145.2000 155.8000 146.0000 160.4000 ;
	    RECT 148.4000 152.2000 149.2000 160.4000 ;
	    RECT 153.2000 153.0000 154.0000 160.4000 ;
	    RECT 161.2000 151.8000 162.0000 160.4000 ;
	    RECT 164.4000 151.8000 165.2000 160.4000 ;
	    RECT 167.6000 151.8000 168.4000 160.4000 ;
	    RECT 170.8000 151.8000 171.6000 160.4000 ;
	    RECT 174.0000 151.8000 174.8000 160.4000 ;
	    RECT 177.2000 153.0000 178.0000 160.4000 ;
	    RECT 183.6000 155.8000 184.4000 160.4000 ;
	    RECT 185.2000 155.8000 186.0000 160.4000 ;
	    RECT 188.4000 155.8000 189.2000 160.4000 ;
	    RECT 191.6000 155.8000 192.4000 160.4000 ;
	    RECT 198.0000 155.8000 198.8000 160.4000 ;
	    RECT 201.2000 155.8000 202.0000 160.4000 ;
	    RECT 209.2000 155.8000 210.0000 160.4000 ;
	    RECT 212.4000 155.8000 213.2000 160.4000 ;
	    RECT 215.6000 155.8000 216.4000 160.4000 ;
	    RECT 218.8000 155.8000 219.6000 160.4000 ;
	    RECT 222.0000 153.0000 222.8000 160.4000 ;
	    RECT 188.4000 151.8000 189.2000 152.4000 ;
	    RECT 191.6000 151.8000 192.6000 152.0000 ;
	    RECT 10.2000 151.2000 37.2000 151.8000 ;
	    RECT 65.2000 151.2000 92.2000 151.8000 ;
	    RECT 100.4000 151.2000 127.4000 151.8000 ;
	    RECT 188.4000 151.2000 215.4000 151.8000 ;
	    RECT 10.2000 151.0000 11.0000 151.2000 ;
	    RECT 91.4000 151.0000 92.2000 151.2000 ;
	    RECT 126.6000 151.0000 127.4000 151.2000 ;
	    RECT 214.6000 151.0000 215.4000 151.2000 ;
	    RECT 153.0000 132.0000 153.8000 132.2000 ;
	    RECT 158.0000 132.0000 158.8000 132.4000 ;
	    RECT 175.6000 132.0000 176.4000 132.6000 ;
	    RECT 153.0000 131.4000 176.4000 132.0000 ;
	    RECT 23.0000 130.8000 23.8000 131.0000 ;
	    RECT 137.8000 130.8000 138.6000 131.0000 ;
	    RECT 216.2000 130.8000 217.0000 131.0000 ;
	    RECT 23.0000 130.2000 50.0000 130.8000 ;
	    RECT 111.6000 130.2000 138.6000 130.8000 ;
	    RECT 190.0000 130.2000 217.0000 130.8000 ;
	    RECT 2.8000 121.6000 3.6000 129.0000 ;
	    RECT 6.0000 121.6000 6.8000 126.2000 ;
	    RECT 10.4000 121.6000 11.2000 130.2000 ;
	    RECT 45.8000 130.0000 46.6000 130.2000 ;
	    RECT 15.6000 121.6000 16.4000 129.8000 ;
	    RECT 49.2000 129.6000 50.0000 130.2000 ;
	    RECT 18.8000 121.6000 19.6000 126.2000 ;
	    RECT 22.0000 121.6000 22.8000 126.2000 ;
	    RECT 25.2000 121.6000 26.0000 126.2000 ;
	    RECT 28.4000 121.6000 29.2000 126.2000 ;
	    RECT 36.4000 121.6000 37.2000 126.2000 ;
	    RECT 39.6000 121.6000 40.4000 126.2000 ;
	    RECT 46.0000 121.6000 46.8000 126.2000 ;
	    RECT 49.2000 121.6000 50.0000 126.2000 ;
	    RECT 52.4000 121.6000 53.2000 126.2000 ;
	    RECT 54.0000 121.6000 54.8000 130.2000 ;
	    RECT 58.2000 121.6000 59.0000 126.2000 ;
	    RECT 62.0000 121.6000 62.8000 129.0000 ;
	    RECT 71.6000 121.6000 72.4000 129.0000 ;
	    RECT 78.0000 121.6000 78.8000 129.0000 ;
	    RECT 82.8000 121.6000 83.6000 129.8000 ;
	    RECT 88.0000 121.6000 88.8000 130.2000 ;
	    RECT 92.4000 121.6000 93.2000 126.2000 ;
	    RECT 94.0000 121.6000 94.8000 130.2000 ;
	    RECT 97.2000 121.6000 98.0000 130.2000 ;
	    RECT 100.4000 121.6000 101.2000 130.2000 ;
	    RECT 103.6000 121.6000 104.4000 130.2000 ;
	    RECT 106.8000 121.6000 107.6000 130.2000 ;
	    RECT 111.6000 129.6000 112.4000 130.2000 ;
	    RECT 114.8000 130.0000 115.8000 130.2000 ;
	    RECT 190.0000 129.6000 190.8000 130.2000 ;
	    RECT 193.4000 130.0000 194.2000 130.2000 ;
	    RECT 108.4000 121.6000 109.2000 126.2000 ;
	    RECT 111.6000 121.6000 112.4000 126.2000 ;
	    RECT 114.8000 121.6000 115.6000 126.2000 ;
	    RECT 121.2000 121.6000 122.0000 126.2000 ;
	    RECT 124.4000 121.6000 125.2000 126.2000 ;
	    RECT 132.4000 121.6000 133.2000 126.2000 ;
	    RECT 135.6000 121.6000 136.4000 126.2000 ;
	    RECT 138.8000 121.6000 139.6000 126.2000 ;
	    RECT 142.0000 121.6000 142.8000 126.2000 ;
	    RECT 143.6000 121.6000 144.4000 126.2000 ;
	    RECT 151.6000 121.6000 152.4000 126.2000 ;
	    RECT 154.8000 121.6000 155.6000 126.2000 ;
	    RECT 158.0000 121.6000 158.8000 126.2000 ;
	    RECT 164.4000 121.6000 165.2000 126.2000 ;
	    RECT 167.6000 121.6000 168.4000 126.2000 ;
	    RECT 175.6000 121.6000 176.4000 126.2000 ;
	    RECT 178.8000 121.6000 179.6000 126.2000 ;
	    RECT 182.0000 121.6000 182.8000 126.2000 ;
	    RECT 185.2000 121.6000 186.0000 126.2000 ;
	    RECT 186.8000 121.6000 187.6000 126.2000 ;
	    RECT 190.0000 121.6000 190.8000 126.2000 ;
	    RECT 193.2000 121.6000 194.0000 126.2000 ;
	    RECT 199.6000 121.6000 200.4000 126.2000 ;
	    RECT 202.8000 121.6000 203.6000 126.2000 ;
	    RECT 210.8000 121.6000 211.6000 126.2000 ;
	    RECT 214.0000 121.6000 214.8000 126.2000 ;
	    RECT 217.2000 121.6000 218.0000 126.2000 ;
	    RECT 220.4000 121.6000 221.2000 126.2000 ;
	    RECT 0.4000 120.4000 226.8000 121.6000 ;
	    RECT 2.8000 113.0000 3.6000 120.4000 ;
	    RECT 7.6000 113.0000 8.4000 120.4000 ;
	    RECT 10.8000 115.8000 11.6000 120.4000 ;
	    RECT 14.0000 115.8000 14.8000 120.4000 ;
	    RECT 18.8000 113.0000 19.6000 120.4000 ;
	    RECT 23.6000 111.8000 24.4000 120.4000 ;
	    RECT 27.8000 115.8000 28.6000 120.4000 ;
	    RECT 31.6000 113.0000 32.4000 120.4000 ;
	    RECT 36.4000 115.8000 37.2000 120.4000 ;
	    RECT 39.6000 115.8000 40.4000 120.4000 ;
	    RECT 42.8000 115.8000 43.6000 120.4000 ;
	    RECT 46.0000 115.8000 46.8000 120.4000 ;
	    RECT 54.0000 115.8000 54.8000 120.4000 ;
	    RECT 57.2000 115.8000 58.0000 120.4000 ;
	    RECT 63.6000 115.8000 64.4000 120.4000 ;
	    RECT 66.8000 115.8000 67.6000 120.4000 ;
	    RECT 70.0000 115.8000 70.8000 120.4000 ;
	    RECT 76.4000 115.8000 77.2000 120.4000 ;
	    RECT 63.4000 111.8000 64.2000 112.0000 ;
	    RECT 66.8000 111.8000 67.6000 112.4000 ;
	    RECT 79.6000 111.8000 80.4000 120.4000 ;
	    RECT 82.8000 111.8000 83.6000 120.4000 ;
	    RECT 86.0000 111.8000 86.8000 120.4000 ;
	    RECT 89.2000 111.8000 90.0000 120.4000 ;
	    RECT 92.4000 111.8000 93.2000 120.4000 ;
	    RECT 94.0000 115.8000 94.8000 120.4000 ;
	    RECT 97.2000 115.8000 98.0000 120.4000 ;
	    RECT 100.4000 115.8000 101.2000 120.4000 ;
	    RECT 106.8000 115.8000 107.6000 120.4000 ;
	    RECT 110.0000 115.8000 110.8000 120.4000 ;
	    RECT 118.0000 115.8000 118.8000 120.4000 ;
	    RECT 121.2000 115.8000 122.0000 120.4000 ;
	    RECT 124.4000 115.8000 125.2000 120.4000 ;
	    RECT 127.6000 115.8000 128.4000 120.4000 ;
	    RECT 129.2000 115.8000 130.0000 120.4000 ;
	    RECT 132.4000 116.2000 133.2000 120.4000 ;
	    RECT 135.6000 115.8000 136.4000 120.4000 ;
	    RECT 97.2000 111.8000 98.0000 112.4000 ;
	    RECT 100.6000 111.8000 101.4000 112.0000 ;
	    RECT 138.8000 111.8000 139.6000 120.4000 ;
	    RECT 145.2000 115.8000 146.0000 120.4000 ;
	    RECT 147.4000 115.8000 148.2000 120.4000 ;
	    RECT 151.6000 111.8000 152.4000 120.4000 ;
	    RECT 153.2000 111.8000 154.0000 120.4000 ;
	    RECT 164.4000 113.0000 165.2000 120.4000 ;
	    RECT 169.2000 111.8000 170.0000 120.4000 ;
	    RECT 173.4000 115.8000 174.2000 120.4000 ;
	    RECT 180.4000 113.0000 181.2000 120.4000 ;
	    RECT 185.2000 115.8000 186.0000 120.4000 ;
	    RECT 188.4000 113.0000 189.2000 120.4000 ;
	    RECT 192.2000 115.8000 193.0000 120.4000 ;
	    RECT 196.4000 111.8000 197.2000 120.4000 ;
	    RECT 198.6000 115.8000 199.4000 120.4000 ;
	    RECT 202.8000 111.8000 203.6000 120.4000 ;
	    RECT 204.4000 115.8000 205.2000 120.4000 ;
	    RECT 207.6000 115.8000 208.4000 120.4000 ;
	    RECT 210.8000 113.0000 211.6000 120.4000 ;
	    RECT 217.2000 115.8000 218.0000 120.4000 ;
	    RECT 220.4000 113.0000 221.2000 120.4000 ;
	    RECT 40.6000 111.2000 67.6000 111.8000 ;
	    RECT 97.2000 111.2000 124.2000 111.8000 ;
	    RECT 40.6000 111.0000 41.4000 111.2000 ;
	    RECT 123.4000 111.0000 124.2000 111.2000 ;
	    RECT 5.4000 90.8000 6.2000 91.0000 ;
	    RECT 72.6000 90.8000 73.4000 91.0000 ;
	    RECT 138.2000 90.8000 139.0000 91.0000 ;
	    RECT 203.4000 90.8000 204.2000 91.0000 ;
	    RECT 5.4000 90.2000 32.4000 90.8000 ;
	    RECT 72.6000 90.2000 99.6000 90.8000 ;
	    RECT 138.2000 90.2000 165.2000 90.8000 ;
	    RECT 28.2000 90.0000 29.0000 90.2000 ;
	    RECT 31.6000 89.6000 32.4000 90.2000 ;
	    RECT 1.2000 81.6000 2.0000 86.2000 ;
	    RECT 4.4000 81.6000 5.2000 86.2000 ;
	    RECT 7.6000 81.6000 8.4000 86.2000 ;
	    RECT 10.8000 81.6000 11.6000 86.2000 ;
	    RECT 18.8000 81.6000 19.6000 86.2000 ;
	    RECT 22.0000 81.6000 22.8000 86.2000 ;
	    RECT 28.4000 81.6000 29.2000 86.2000 ;
	    RECT 31.6000 81.6000 32.4000 86.2000 ;
	    RECT 34.8000 81.6000 35.6000 86.2000 ;
	    RECT 38.0000 81.6000 38.8000 89.0000 ;
	    RECT 41.8000 81.6000 42.6000 86.2000 ;
	    RECT 46.0000 81.6000 46.8000 90.2000 ;
	    RECT 95.4000 90.0000 96.2000 90.2000 ;
	    RECT 98.8000 89.6000 99.6000 90.2000 ;
	    RECT 161.0000 90.0000 161.8000 90.2000 ;
	    RECT 164.4000 89.6000 165.2000 90.2000 ;
	    RECT 177.2000 90.2000 204.2000 90.8000 ;
	    RECT 177.2000 89.6000 178.0000 90.2000 ;
	    RECT 180.4000 90.0000 181.4000 90.2000 ;
	    RECT 49.2000 81.6000 50.2000 88.8000 ;
	    RECT 55.4000 82.2000 56.4000 88.8000 ;
	    RECT 55.4000 81.6000 56.2000 82.2000 ;
	    RECT 60.4000 81.6000 61.2000 89.0000 ;
	    RECT 68.4000 81.6000 69.2000 86.2000 ;
	    RECT 71.6000 81.6000 72.4000 86.2000 ;
	    RECT 74.8000 81.6000 75.6000 86.2000 ;
	    RECT 78.0000 81.6000 78.8000 86.2000 ;
	    RECT 86.0000 81.6000 86.8000 86.2000 ;
	    RECT 89.2000 81.6000 90.0000 86.2000 ;
	    RECT 95.6000 81.6000 96.4000 86.2000 ;
	    RECT 98.8000 81.6000 99.6000 86.2000 ;
	    RECT 102.0000 81.6000 102.8000 86.2000 ;
	    RECT 105.2000 81.6000 106.0000 89.0000 ;
	    RECT 110.0000 81.6000 110.8000 89.0000 ;
	    RECT 114.8000 81.6000 115.6000 89.0000 ;
	    RECT 119.6000 81.6000 120.4000 85.8000 ;
	    RECT 122.8000 81.6000 123.6000 86.2000 ;
	    RECT 124.4000 81.6000 125.2000 86.2000 ;
	    RECT 127.6000 81.6000 128.4000 85.8000 ;
	    RECT 132.4000 81.6000 133.2000 86.2000 ;
	    RECT 134.0000 81.6000 134.8000 86.2000 ;
	    RECT 137.2000 81.6000 138.0000 86.2000 ;
	    RECT 140.4000 81.6000 141.2000 86.2000 ;
	    RECT 143.6000 81.6000 144.4000 86.2000 ;
	    RECT 151.6000 81.6000 152.4000 86.2000 ;
	    RECT 154.8000 81.6000 155.6000 86.2000 ;
	    RECT 161.2000 81.6000 162.0000 86.2000 ;
	    RECT 164.4000 81.6000 165.2000 86.2000 ;
	    RECT 167.6000 81.6000 168.4000 86.2000 ;
	    RECT 174.0000 81.6000 174.8000 86.2000 ;
	    RECT 177.2000 81.6000 178.0000 86.2000 ;
	    RECT 180.4000 81.6000 181.2000 86.2000 ;
	    RECT 186.8000 81.6000 187.6000 86.2000 ;
	    RECT 190.0000 81.6000 190.8000 86.2000 ;
	    RECT 198.0000 81.6000 198.8000 86.2000 ;
	    RECT 201.2000 81.6000 202.0000 86.2000 ;
	    RECT 204.4000 81.6000 205.2000 86.2000 ;
	    RECT 207.6000 81.6000 208.4000 86.2000 ;
	    RECT 209.2000 81.6000 210.0000 86.2000 ;
	    RECT 212.4000 81.6000 213.2000 86.2000 ;
	    RECT 214.0000 81.6000 214.8000 90.2000 ;
	    RECT 218.2000 81.6000 219.0000 86.2000 ;
	    RECT 220.4000 81.6000 221.2000 86.2000 ;
	    RECT 223.6000 81.6000 224.4000 85.8000 ;
	    RECT 0.4000 80.4000 226.8000 81.6000 ;
	    RECT 1.2000 75.8000 2.0000 80.4000 ;
	    RECT 4.4000 75.8000 5.2000 80.4000 ;
	    RECT 7.6000 75.8000 8.4000 80.4000 ;
	    RECT 10.8000 75.8000 11.6000 80.4000 ;
	    RECT 18.8000 75.8000 19.6000 80.4000 ;
	    RECT 22.0000 75.8000 22.8000 80.4000 ;
	    RECT 28.4000 75.8000 29.2000 80.4000 ;
	    RECT 31.6000 75.8000 32.4000 80.4000 ;
	    RECT 34.8000 75.8000 35.6000 80.4000 ;
	    RECT 28.2000 71.8000 29.0000 72.0000 ;
	    RECT 31.6000 71.8000 32.4000 72.4000 ;
	    RECT 36.4000 71.8000 37.2000 80.4000 ;
	    RECT 40.6000 75.8000 41.4000 80.4000 ;
	    RECT 43.4000 75.8000 44.2000 80.4000 ;
	    RECT 47.6000 71.8000 48.4000 80.4000 ;
	    RECT 50.8000 73.0000 51.6000 80.4000 ;
	    RECT 55.6000 71.8000 56.4000 80.4000 ;
	    RECT 59.8000 75.8000 60.6000 80.4000 ;
	    RECT 66.8000 75.8000 67.6000 80.4000 ;
	    RECT 73.2000 71.8000 74.0000 80.4000 ;
	    RECT 75.4000 75.8000 76.2000 80.4000 ;
	    RECT 79.6000 71.8000 80.4000 80.4000 ;
	    RECT 81.2000 75.8000 82.0000 80.4000 ;
	    RECT 84.4000 75.8000 85.2000 80.4000 ;
	    RECT 87.6000 75.8000 88.4000 80.4000 ;
	    RECT 94.0000 75.8000 94.8000 80.4000 ;
	    RECT 97.2000 75.8000 98.0000 80.4000 ;
	    RECT 105.2000 75.8000 106.0000 80.4000 ;
	    RECT 108.4000 75.8000 109.2000 80.4000 ;
	    RECT 111.6000 75.8000 112.4000 80.4000 ;
	    RECT 114.8000 75.8000 115.6000 80.4000 ;
	    RECT 116.4000 75.8000 117.2000 80.4000 ;
	    RECT 121.2000 75.8000 122.0000 80.4000 ;
	    RECT 124.4000 73.0000 125.2000 80.4000 ;
	    RECT 132.4000 73.8000 133.2000 80.4000 ;
	    RECT 148.4000 75.8000 149.2000 80.4000 ;
	    RECT 151.6000 75.8000 152.4000 80.4000 ;
	    RECT 154.8000 75.8000 155.6000 80.4000 ;
	    RECT 161.2000 75.8000 162.0000 80.4000 ;
	    RECT 164.4000 75.8000 165.2000 80.4000 ;
	    RECT 172.4000 75.8000 173.2000 80.4000 ;
	    RECT 175.6000 75.8000 176.4000 80.4000 ;
	    RECT 178.8000 75.8000 179.6000 80.4000 ;
	    RECT 182.0000 75.8000 182.8000 80.4000 ;
	    RECT 84.4000 71.8000 85.2000 72.4000 ;
	    RECT 87.6000 71.8000 88.6000 72.0000 ;
	    RECT 151.6000 71.8000 152.4000 72.4000 ;
	    RECT 155.0000 71.8000 155.8000 72.0000 ;
	    RECT 183.6000 71.8000 184.4000 80.4000 ;
	    RECT 187.8000 75.8000 188.6000 80.4000 ;
	    RECT 190.0000 71.8000 190.8000 80.4000 ;
	    RECT 194.2000 75.8000 195.0000 80.4000 ;
	    RECT 199.6000 73.0000 200.4000 80.4000 ;
	    RECT 203.4000 75.8000 204.2000 80.4000 ;
	    RECT 207.6000 71.8000 208.4000 80.4000 ;
	    RECT 209.2000 75.8000 210.0000 80.4000 ;
	    RECT 212.4000 76.2000 213.2000 80.4000 ;
	    RECT 215.6000 71.8000 216.4000 80.4000 ;
	    RECT 219.8000 75.8000 220.6000 80.4000 ;
	    RECT 225.2000 71.8000 226.0000 80.4000 ;
	    RECT 5.4000 71.2000 32.4000 71.8000 ;
	    RECT 84.4000 71.2000 111.4000 71.8000 ;
	    RECT 151.6000 71.2000 178.6000 71.8000 ;
	    RECT 5.4000 71.0000 6.2000 71.2000 ;
	    RECT 110.6000 71.0000 111.4000 71.2000 ;
	    RECT 177.8000 71.0000 178.6000 71.2000 ;
	    RECT 128.6000 50.8000 129.4000 51.0000 ;
	    RECT 128.6000 50.2000 155.6000 50.8000 ;
	    RECT 2.8000 41.6000 3.6000 49.0000 ;
	    RECT 7.6000 41.6000 8.4000 49.0000 ;
	    RECT 12.0000 41.6000 12.8000 50.2000 ;
	    RECT 17.2000 41.6000 18.0000 49.8000 ;
	    RECT 22.0000 41.6000 22.8000 46.2000 ;
	    RECT 25.2000 41.6000 26.0000 49.0000 ;
	    RECT 31.6000 41.6000 32.4000 49.0000 ;
	    RECT 38.0000 41.6000 38.8000 46.2000 ;
	    RECT 41.2000 41.6000 42.2000 48.8000 ;
	    RECT 47.4000 42.2000 48.4000 48.8000 ;
	    RECT 47.4000 41.6000 48.2000 42.2000 ;
	    RECT 52.4000 41.6000 53.2000 49.8000 ;
	    RECT 57.6000 41.6000 58.4000 50.2000 ;
	    RECT 62.0000 41.6000 62.8000 49.0000 ;
	    RECT 71.6000 41.6000 72.4000 46.2000 ;
	    RECT 73.2000 41.6000 74.0000 50.2000 ;
	    RECT 76.4000 41.6000 77.2000 50.2000 ;
	    RECT 79.6000 41.6000 80.4000 50.2000 ;
	    RECT 82.8000 41.6000 83.6000 50.2000 ;
	    RECT 86.0000 41.6000 86.8000 50.2000 ;
	    RECT 87.6000 41.6000 88.4000 50.2000 ;
	    RECT 90.8000 41.6000 91.6000 50.2000 ;
	    RECT 94.0000 41.6000 94.8000 50.2000 ;
	    RECT 97.2000 41.6000 98.0000 50.2000 ;
	    RECT 100.4000 41.6000 101.2000 50.2000 ;
	    RECT 102.0000 41.6000 102.8000 50.2000 ;
	    RECT 151.4000 50.0000 152.2000 50.2000 ;
	    RECT 154.8000 49.6000 155.6000 50.2000 ;
	    RECT 106.8000 41.6000 107.6000 46.2000 ;
	    RECT 110.0000 41.6000 110.8000 46.2000 ;
	    RECT 111.6000 41.6000 112.4000 46.2000 ;
	    RECT 114.8000 41.6000 115.6000 45.8000 ;
	    RECT 119.6000 41.6000 120.4000 45.8000 ;
	    RECT 122.8000 41.6000 123.6000 46.2000 ;
	    RECT 124.4000 41.6000 125.2000 46.2000 ;
	    RECT 127.6000 41.6000 128.4000 46.2000 ;
	    RECT 130.8000 41.6000 131.6000 46.2000 ;
	    RECT 134.0000 41.6000 134.8000 46.2000 ;
	    RECT 142.0000 41.6000 142.8000 46.2000 ;
	    RECT 145.2000 41.6000 146.0000 46.2000 ;
	    RECT 151.6000 41.6000 152.4000 46.2000 ;
	    RECT 154.8000 41.6000 155.6000 46.2000 ;
	    RECT 158.0000 41.6000 158.8000 46.2000 ;
	    RECT 164.4000 41.6000 165.2000 50.2000 ;
	    RECT 168.6000 41.6000 169.4000 46.2000 ;
	    RECT 170.8000 41.6000 171.6000 46.2000 ;
	    RECT 174.0000 41.6000 174.8000 49.8000 ;
	    RECT 177.8000 41.6000 178.6000 46.2000 ;
	    RECT 182.0000 41.6000 182.8000 50.2000 ;
	    RECT 186.8000 41.6000 187.6000 50.2000 ;
	    RECT 190.0000 42.2000 191.0000 48.8000 ;
	    RECT 190.2000 41.6000 191.0000 42.2000 ;
	    RECT 196.2000 41.6000 197.2000 48.8000 ;
	    RECT 200.2000 41.6000 201.0000 46.2000 ;
	    RECT 204.4000 41.6000 205.2000 50.2000 ;
	    RECT 207.6000 41.6000 208.4000 49.0000 ;
	    RECT 210.8000 41.6000 211.6000 46.2000 ;
	    RECT 214.0000 41.6000 214.8000 50.2000 ;
	    RECT 218.8000 41.6000 219.6000 46.2000 ;
	    RECT 222.0000 41.6000 222.8000 46.2000 ;
	    RECT 0.4000 40.4000 226.8000 41.6000 ;
	    RECT 1.2000 35.8000 2.0000 40.4000 ;
	    RECT 4.4000 35.8000 5.2000 40.4000 ;
	    RECT 7.6000 35.8000 8.4000 40.4000 ;
	    RECT 10.8000 35.8000 11.6000 40.4000 ;
	    RECT 14.0000 35.8000 14.8000 40.4000 ;
	    RECT 22.0000 35.8000 22.8000 40.4000 ;
	    RECT 25.2000 35.8000 26.0000 40.4000 ;
	    RECT 31.6000 35.8000 32.4000 40.4000 ;
	    RECT 34.8000 35.8000 35.6000 40.4000 ;
	    RECT 38.0000 35.8000 38.8000 40.4000 ;
	    RECT 39.6000 35.8000 40.4000 40.4000 ;
	    RECT 42.8000 35.8000 43.6000 40.4000 ;
	    RECT 46.0000 35.8000 46.8000 40.4000 ;
	    RECT 52.4000 35.8000 53.2000 40.4000 ;
	    RECT 55.6000 35.8000 56.4000 40.4000 ;
	    RECT 63.6000 35.8000 64.4000 40.4000 ;
	    RECT 66.8000 35.8000 67.6000 40.4000 ;
	    RECT 70.0000 35.8000 70.8000 40.4000 ;
	    RECT 73.2000 35.8000 74.0000 40.4000 ;
	    RECT 79.6000 35.8000 80.4000 40.4000 ;
	    RECT 82.8000 35.8000 83.6000 40.4000 ;
	    RECT 85.0000 35.8000 85.8000 40.4000 ;
	    RECT 31.4000 31.8000 32.2000 32.0000 ;
	    RECT 34.8000 31.8000 35.6000 32.4000 ;
	    RECT 8.6000 31.2000 35.6000 31.8000 ;
	    RECT 42.8000 31.8000 43.6000 32.4000 ;
	    RECT 46.0000 31.8000 47.0000 32.0000 ;
	    RECT 89.2000 31.8000 90.0000 40.4000 ;
	    RECT 90.8000 31.8000 91.6000 40.4000 ;
	    RECT 95.0000 35.8000 95.8000 40.4000 ;
	    RECT 97.2000 35.8000 98.0000 40.4000 ;
	    RECT 100.4000 35.8000 101.2000 40.4000 ;
	    RECT 103.6000 36.2000 104.4000 40.4000 ;
	    RECT 108.4000 36.2000 109.2000 40.4000 ;
	    RECT 111.6000 35.8000 112.4000 40.4000 ;
	    RECT 114.8000 32.2000 115.6000 40.4000 ;
	    RECT 118.0000 35.8000 118.8000 40.4000 ;
	    RECT 119.6000 31.8000 120.4000 40.4000 ;
	    RECT 124.4000 35.8000 125.2000 40.4000 ;
	    RECT 127.6000 35.8000 128.4000 40.4000 ;
	    RECT 130.8000 35.8000 131.6000 40.4000 ;
	    RECT 134.0000 35.8000 134.8000 40.4000 ;
	    RECT 142.0000 35.8000 142.8000 40.4000 ;
	    RECT 145.2000 35.8000 146.0000 40.4000 ;
	    RECT 151.6000 35.8000 152.4000 40.4000 ;
	    RECT 154.8000 35.8000 155.6000 40.4000 ;
	    RECT 158.0000 35.8000 158.8000 40.4000 ;
	    RECT 164.4000 35.8000 165.2000 40.4000 ;
	    RECT 167.6000 35.8000 168.4000 40.4000 ;
	    RECT 170.8000 35.8000 171.6000 40.4000 ;
	    RECT 151.4000 31.8000 152.2000 32.0000 ;
	    RECT 154.8000 31.8000 155.6000 32.4000 ;
	    RECT 175.6000 31.8000 176.4000 40.4000 ;
	    RECT 177.2000 35.8000 178.0000 40.4000 ;
	    RECT 180.4000 31.8000 181.2000 40.4000 ;
	    RECT 184.6000 35.8000 185.4000 40.4000 ;
	    RECT 186.8000 35.8000 187.6000 40.4000 ;
	    RECT 190.0000 35.8000 190.8000 40.4000 ;
	    RECT 191.6000 35.8000 192.4000 40.4000 ;
	    RECT 194.8000 36.2000 195.6000 40.4000 ;
	    RECT 198.6000 35.8000 199.4000 40.4000 ;
	    RECT 202.8000 31.8000 203.6000 40.4000 ;
	    RECT 204.4000 35.8000 205.2000 40.4000 ;
	    RECT 208.2000 35.8000 209.0000 40.4000 ;
	    RECT 212.4000 31.8000 213.2000 40.4000 ;
	    RECT 214.0000 35.8000 214.8000 40.4000 ;
	    RECT 217.2000 36.2000 218.0000 40.4000 ;
	    RECT 220.4000 31.8000 221.2000 40.4000 ;
	    RECT 42.8000 31.2000 69.8000 31.8000 ;
	    RECT 8.6000 31.0000 9.4000 31.2000 ;
	    RECT 69.0000 31.0000 69.8000 31.2000 ;
	    RECT 128.6000 31.2000 155.6000 31.8000 ;
	    RECT 128.6000 31.0000 129.4000 31.2000 ;
	    RECT 10.2000 10.8000 11.0000 11.0000 ;
	    RECT 70.6000 10.8000 71.4000 11.0000 ;
	    RECT 10.2000 10.2000 37.2000 10.8000 ;
	    RECT 33.0000 10.0000 33.8000 10.2000 ;
	    RECT 36.4000 9.6000 37.2000 10.2000 ;
	    RECT 44.4000 10.2000 71.4000 10.8000 ;
	    RECT 95.0000 10.8000 95.8000 11.0000 ;
	    RECT 173.4000 10.8000 174.2000 11.0000 ;
	    RECT 95.0000 10.2000 122.0000 10.8000 ;
	    RECT 173.4000 10.2000 200.4000 10.8000 ;
	    RECT 44.4000 9.6000 45.2000 10.2000 ;
	    RECT 47.8000 10.0000 48.6000 10.2000 ;
	    RECT 117.8000 10.0000 118.6000 10.2000 ;
	    RECT 121.2000 9.6000 122.0000 10.2000 ;
	    RECT 2.8000 1.6000 3.6000 9.0000 ;
	    RECT 6.0000 1.6000 6.8000 6.2000 ;
	    RECT 9.2000 1.6000 10.0000 6.2000 ;
	    RECT 12.4000 1.6000 13.2000 6.2000 ;
	    RECT 15.6000 1.6000 16.4000 6.2000 ;
	    RECT 23.6000 1.6000 24.4000 6.2000 ;
	    RECT 26.8000 1.6000 27.6000 6.2000 ;
	    RECT 33.2000 1.6000 34.0000 6.2000 ;
	    RECT 36.4000 1.6000 37.2000 6.2000 ;
	    RECT 39.6000 1.6000 40.4000 6.2000 ;
	    RECT 41.2000 1.6000 42.0000 6.2000 ;
	    RECT 44.4000 1.6000 45.2000 6.2000 ;
	    RECT 47.6000 1.6000 48.4000 6.2000 ;
	    RECT 54.0000 1.6000 54.8000 6.2000 ;
	    RECT 57.2000 1.6000 58.0000 6.2000 ;
	    RECT 65.2000 1.6000 66.0000 6.2000 ;
	    RECT 68.4000 1.6000 69.2000 6.2000 ;
	    RECT 71.6000 1.6000 72.4000 6.2000 ;
	    RECT 74.8000 1.6000 75.6000 6.2000 ;
	    RECT 82.8000 1.6000 83.6000 9.0000 ;
	    RECT 87.6000 1.6000 88.4000 9.0000 ;
	    RECT 90.8000 1.6000 91.6000 6.2000 ;
	    RECT 94.0000 1.6000 94.8000 6.2000 ;
	    RECT 97.2000 1.6000 98.0000 6.2000 ;
	    RECT 100.4000 1.6000 101.2000 6.2000 ;
	    RECT 108.4000 1.6000 109.2000 6.2000 ;
	    RECT 111.6000 1.6000 112.4000 6.2000 ;
	    RECT 118.0000 1.6000 118.8000 6.2000 ;
	    RECT 121.2000 1.6000 122.0000 6.2000 ;
	    RECT 124.4000 1.6000 125.2000 6.2000 ;
	    RECT 127.6000 1.6000 128.4000 9.0000 ;
	    RECT 132.4000 1.6000 133.2000 9.0000 ;
	    RECT 135.6000 1.6000 136.4000 10.2000 ;
	    RECT 140.4000 1.6000 141.2000 6.2000 ;
	    RECT 143.6000 1.6000 144.4000 9.8000 ;
	    RECT 146.8000 1.6000 147.6000 10.2000 ;
	    RECT 151.0000 1.6000 151.8000 6.2000 ;
	    RECT 153.8000 1.6000 154.6000 6.2000 ;
	    RECT 158.0000 1.6000 158.8000 10.2000 ;
	    RECT 196.2000 10.0000 197.0000 10.2000 ;
	    RECT 199.6000 9.6000 200.4000 10.2000 ;
	    RECT 166.0000 1.6000 166.8000 9.0000 ;
	    RECT 169.2000 1.6000 170.0000 6.2000 ;
	    RECT 172.4000 1.6000 173.2000 6.2000 ;
	    RECT 175.6000 1.6000 176.4000 6.2000 ;
	    RECT 178.8000 1.6000 179.6000 6.2000 ;
	    RECT 186.8000 1.6000 187.6000 6.2000 ;
	    RECT 190.0000 1.6000 190.8000 6.2000 ;
	    RECT 196.4000 1.6000 197.2000 6.2000 ;
	    RECT 199.6000 1.6000 200.4000 6.2000 ;
	    RECT 202.8000 1.6000 203.6000 6.2000 ;
	    RECT 204.4000 1.6000 205.2000 10.2000 ;
	    RECT 208.6000 1.6000 209.4000 6.2000 ;
	    RECT 212.4000 1.6000 213.2000 6.2000 ;
	    RECT 215.6000 1.6000 216.4000 6.2000 ;
	    RECT 218.8000 1.6000 219.6000 6.2000 ;
	    RECT 222.0000 1.6000 222.8000 9.0000 ;
	    RECT 0.4000 0.4000 226.8000 1.6000 ;
         LAYER metal2 ;
	    RECT 63.2000 200.6000 68.0000 201.4000 ;
	    RECT 36.4000 197.6000 37.2000 198.4000 ;
	    RECT 81.2000 197.6000 82.0000 198.4000 ;
	    RECT 196.4000 197.6000 197.2000 198.4000 ;
	    RECT 36.5000 192.4000 37.1000 197.6000 ;
	    RECT 81.3000 192.4000 81.9000 197.6000 ;
	    RECT 121.2000 195.8000 122.0000 196.6000 ;
	    RECT 36.4000 191.6000 37.2000 192.4000 ;
	    RECT 81.2000 191.6000 82.0000 192.4000 ;
	    RECT 121.3000 192.0000 121.9000 195.8000 ;
	    RECT 196.5000 192.4000 197.1000 197.6000 ;
	    RECT 121.2000 191.2000 122.0000 192.0000 ;
	    RECT 196.4000 191.6000 197.2000 192.4000 ;
	    RECT 46.0000 170.0000 46.8000 170.8000 ;
	    RECT 114.8000 170.0000 115.6000 170.8000 ;
	    RECT 46.1000 164.4000 46.7000 170.0000 ;
	    RECT 114.9000 166.2000 115.5000 170.0000 ;
	    RECT 186.8000 169.6000 187.6000 170.4000 ;
	    RECT 194.8000 169.6000 195.6000 170.4000 ;
	    RECT 114.8000 165.4000 115.6000 166.2000 ;
	    RECT 186.9000 164.4000 187.5000 169.6000 ;
	    RECT 194.9000 164.4000 195.5000 169.6000 ;
	    RECT 46.0000 163.6000 46.8000 164.4000 ;
	    RECT 186.8000 163.6000 187.6000 164.4000 ;
	    RECT 194.8000 163.6000 195.6000 164.4000 ;
	    RECT 63.2000 160.6000 68.0000 161.4000 ;
	    RECT 36.4000 157.6000 37.2000 158.4000 ;
	    RECT 65.2000 157.6000 66.0000 158.4000 ;
	    RECT 36.5000 152.4000 37.1000 157.6000 ;
	    RECT 65.3000 152.4000 65.9000 157.6000 ;
	    RECT 103.6000 155.8000 104.4000 156.6000 ;
	    RECT 191.6000 155.8000 192.4000 156.6000 ;
	    RECT 36.4000 151.6000 37.2000 152.4000 ;
	    RECT 65.2000 151.6000 66.0000 152.4000 ;
	    RECT 103.7000 152.0000 104.3000 155.8000 ;
	    RECT 191.7000 152.0000 192.3000 155.8000 ;
	    RECT 103.6000 151.2000 104.4000 152.0000 ;
	    RECT 191.6000 151.2000 192.4000 152.0000 ;
	    RECT 175.6000 131.6000 176.4000 132.4000 ;
	    RECT 49.2000 129.6000 50.0000 130.4000 ;
	    RECT 114.8000 130.0000 115.6000 130.8000 ;
	    RECT 49.3000 124.4000 49.9000 129.6000 ;
	    RECT 114.9000 124.4000 115.5000 130.0000 ;
	    RECT 175.7000 126.2000 176.3000 131.6000 ;
	    RECT 190.0000 129.6000 190.8000 130.4000 ;
	    RECT 175.6000 125.4000 176.4000 126.2000 ;
	    RECT 190.1000 124.4000 190.7000 129.6000 ;
	    RECT 49.2000 123.6000 50.0000 124.4000 ;
	    RECT 114.8000 123.6000 115.6000 124.4000 ;
	    RECT 190.0000 123.6000 190.8000 124.4000 ;
	    RECT 63.2000 120.6000 68.0000 121.4000 ;
	    RECT 66.8000 117.6000 67.6000 118.4000 ;
	    RECT 97.2000 117.6000 98.0000 118.4000 ;
	    RECT 66.9000 112.4000 67.5000 117.6000 ;
	    RECT 97.3000 112.4000 97.9000 117.6000 ;
	    RECT 66.8000 111.6000 67.6000 112.4000 ;
	    RECT 97.2000 111.6000 98.0000 112.4000 ;
	    RECT 31.6000 89.6000 32.4000 90.4000 ;
	    RECT 98.8000 89.6000 99.6000 90.4000 ;
	    RECT 164.4000 89.6000 165.2000 90.4000 ;
	    RECT 180.4000 90.0000 181.2000 90.8000 ;
	    RECT 31.7000 84.4000 32.3000 89.6000 ;
	    RECT 98.9000 84.4000 99.5000 89.6000 ;
	    RECT 164.5000 84.4000 165.1000 89.6000 ;
	    RECT 180.5000 86.2000 181.1000 90.0000 ;
	    RECT 180.4000 85.4000 181.2000 86.2000 ;
	    RECT 31.6000 83.6000 32.4000 84.4000 ;
	    RECT 98.8000 83.6000 99.6000 84.4000 ;
	    RECT 164.4000 83.6000 165.2000 84.4000 ;
	    RECT 63.2000 80.6000 68.0000 81.4000 ;
	    RECT 31.6000 77.6000 32.4000 78.4000 ;
	    RECT 151.6000 77.6000 152.4000 78.4000 ;
	    RECT 31.7000 72.4000 32.3000 77.6000 ;
	    RECT 87.6000 75.8000 88.4000 76.6000 ;
	    RECT 31.6000 71.6000 32.4000 72.4000 ;
	    RECT 87.7000 72.0000 88.3000 75.8000 ;
	    RECT 151.7000 72.4000 152.3000 77.6000 ;
	    RECT 87.6000 71.2000 88.4000 72.0000 ;
	    RECT 151.6000 71.6000 152.4000 72.4000 ;
	    RECT 154.8000 49.6000 155.6000 50.4000 ;
	    RECT 154.9000 44.4000 155.5000 49.6000 ;
	    RECT 154.8000 43.6000 155.6000 44.4000 ;
	    RECT 63.2000 40.6000 68.0000 41.4000 ;
	    RECT 34.8000 37.6000 35.6000 38.4000 ;
	    RECT 154.8000 37.6000 155.6000 38.4000 ;
	    RECT 34.9000 32.4000 35.5000 37.6000 ;
	    RECT 46.0000 35.8000 46.8000 36.6000 ;
	    RECT 34.8000 31.6000 35.6000 32.4000 ;
	    RECT 46.1000 32.0000 46.7000 35.8000 ;
	    RECT 154.9000 32.4000 155.5000 37.6000 ;
	    RECT 46.0000 31.2000 46.8000 32.0000 ;
	    RECT 154.8000 31.6000 155.6000 32.4000 ;
	    RECT 36.4000 9.6000 37.2000 10.4000 ;
	    RECT 44.4000 9.6000 45.2000 10.4000 ;
	    RECT 121.2000 9.6000 122.0000 10.4000 ;
	    RECT 199.6000 9.6000 200.4000 10.4000 ;
	    RECT 36.5000 4.4000 37.1000 9.6000 ;
	    RECT 44.5000 4.4000 45.1000 9.6000 ;
	    RECT 121.3000 4.4000 121.9000 9.6000 ;
	    RECT 199.7000 4.4000 200.3000 9.6000 ;
	    RECT 36.4000 3.6000 37.2000 4.4000 ;
	    RECT 44.4000 3.6000 45.2000 4.4000 ;
	    RECT 121.2000 3.6000 122.0000 4.4000 ;
	    RECT 199.6000 3.6000 200.4000 4.4000 ;
	    RECT 63.2000 0.6000 68.0000 1.4000 ;
         LAYER metal3 ;
	    RECT 63.2000 200.4000 68.0000 201.6000 ;
	    RECT 63.2000 160.4000 68.0000 161.6000 ;
	    RECT 63.2000 120.4000 68.0000 121.6000 ;
	    RECT 63.2000 80.4000 68.0000 81.6000 ;
	    RECT 63.2000 40.4000 68.0000 41.6000 ;
	    RECT 63.2000 0.4000 68.0000 1.6000 ;
         LAYER metal4 ;
	    RECT 63.2000 -4.0000 68.0000 204.0000 ;
      END
   END vdd
   PIN gnd
      PORT
         LAYER metal1 ;
	    RECT 2.8000 181.6000 3.6000 186.2000 ;
	    RECT 6.0000 181.6000 6.8000 184.2000 ;
	    RECT 12.4000 181.6000 13.2000 186.2000 ;
	    RECT 23.6000 181.6000 24.4000 184.2000 ;
	    RECT 26.8000 181.6000 27.6000 184.2000 ;
	    RECT 36.4000 181.6000 37.2000 186.2000 ;
	    RECT 42.8000 181.6000 43.6000 186.2000 ;
	    RECT 50.8000 181.6000 51.6000 184.2000 ;
	    RECT 57.2000 181.6000 58.0000 186.2000 ;
	    RECT 68.4000 181.6000 69.2000 184.2000 ;
	    RECT 71.6000 181.6000 72.4000 184.2000 ;
	    RECT 81.2000 181.6000 82.0000 186.2000 ;
	    RECT 87.6000 181.6000 88.4000 186.2000 ;
	    RECT 92.4000 181.6000 93.2000 186.2000 ;
	    RECT 97.2000 181.6000 98.0000 186.2000 ;
	    RECT 100.4000 181.6000 101.2000 184.2000 ;
	    RECT 104.2000 181.6000 105.0000 186.2000 ;
	    RECT 108.4000 181.6000 109.2000 184.2000 ;
	    RECT 110.0000 181.6000 110.8000 184.2000 ;
	    RECT 113.2000 181.6000 114.0000 184.2000 ;
	    RECT 118.0000 181.6000 118.8000 186.2000 ;
	    RECT 127.6000 181.6000 128.4000 184.2000 ;
	    RECT 130.8000 181.6000 131.6000 184.2000 ;
	    RECT 142.0000 181.6000 142.8000 186.2000 ;
	    RECT 148.4000 181.6000 149.2000 184.2000 ;
	    RECT 150.0000 181.6000 150.8000 188.2000 ;
	    RECT 162.8000 181.6000 163.6000 186.2000 ;
	    RECT 166.0000 181.6000 166.8000 184.2000 ;
	    RECT 172.4000 181.6000 173.2000 186.2000 ;
	    RECT 183.6000 181.6000 184.4000 184.2000 ;
	    RECT 186.8000 181.6000 187.6000 184.2000 ;
	    RECT 196.4000 181.6000 197.2000 186.2000 ;
	    RECT 201.2000 181.6000 202.0000 184.2000 ;
	    RECT 204.4000 181.6000 205.2000 184.2000 ;
	    RECT 206.0000 181.6000 206.8000 184.2000 ;
	    RECT 210.2000 181.6000 211.0000 186.2000 ;
	    RECT 214.0000 181.6000 214.8000 184.2000 ;
	    RECT 217.2000 181.6000 218.0000 186.2000 ;
	    RECT 222.0000 181.6000 222.8000 184.2000 ;
	    RECT 0.4000 180.4000 226.8000 181.6000 ;
	    RECT 2.8000 175.8000 3.6000 180.4000 ;
	    RECT 6.0000 177.8000 6.8000 180.4000 ;
	    RECT 10.4000 175.0000 11.2000 180.4000 ;
	    RECT 15.6000 175.4000 16.4000 180.4000 ;
	    RECT 18.8000 177.8000 19.6000 180.4000 ;
	    RECT 25.2000 175.8000 26.0000 180.4000 ;
	    RECT 36.4000 177.8000 37.2000 180.4000 ;
	    RECT 39.6000 177.8000 40.4000 180.4000 ;
	    RECT 49.2000 175.8000 50.0000 180.4000 ;
	    RECT 54.0000 177.8000 54.8000 180.4000 ;
	    RECT 57.2000 177.8000 58.0000 180.4000 ;
	    RECT 66.4000 175.0000 67.2000 180.4000 ;
	    RECT 71.6000 175.4000 72.4000 180.4000 ;
	    RECT 75.4000 175.8000 76.2000 180.4000 ;
	    RECT 79.6000 177.8000 80.4000 180.4000 ;
	    RECT 82.8000 176.6000 83.6000 180.4000 ;
	    RECT 87.6000 177.8000 88.4000 180.4000 ;
	    RECT 94.0000 175.8000 94.8000 180.4000 ;
	    RECT 105.2000 177.8000 106.0000 180.4000 ;
	    RECT 108.4000 177.8000 109.2000 180.4000 ;
	    RECT 118.0000 175.8000 118.8000 180.4000 ;
	    RECT 124.4000 175.8000 125.2000 180.4000 ;
	    RECT 129.2000 175.4000 130.0000 180.4000 ;
	    RECT 134.4000 175.0000 135.2000 180.4000 ;
	    RECT 138.8000 177.8000 139.6000 180.4000 ;
	    RECT 142.0000 177.8000 142.8000 180.4000 ;
	    RECT 143.6000 177.8000 144.4000 180.4000 ;
	    RECT 146.8000 177.8000 147.6000 180.4000 ;
	    RECT 150.0000 177.8000 150.8000 180.4000 ;
	    RECT 156.4000 177.8000 157.2000 180.4000 ;
	    RECT 162.8000 175.8000 163.6000 180.4000 ;
	    RECT 174.0000 177.8000 174.8000 180.4000 ;
	    RECT 177.2000 177.8000 178.0000 180.4000 ;
	    RECT 186.8000 175.8000 187.6000 180.4000 ;
	    RECT 194.8000 175.8000 195.6000 180.4000 ;
	    RECT 204.4000 177.8000 205.2000 180.4000 ;
	    RECT 207.6000 177.8000 208.4000 180.4000 ;
	    RECT 218.8000 175.8000 219.6000 180.4000 ;
	    RECT 225.2000 177.8000 226.0000 180.4000 ;
	    RECT 2.8000 141.6000 3.6000 146.2000 ;
	    RECT 6.0000 141.6000 6.8000 144.2000 ;
	    RECT 12.4000 141.6000 13.2000 146.2000 ;
	    RECT 23.6000 141.6000 24.4000 144.2000 ;
	    RECT 26.8000 141.6000 27.6000 144.2000 ;
	    RECT 36.4000 141.6000 37.2000 146.2000 ;
	    RECT 44.4000 141.6000 45.2000 145.4000 ;
	    RECT 47.6000 141.6000 48.4000 144.2000 ;
	    RECT 51.8000 141.6000 52.6000 146.2000 ;
	    RECT 54.0000 141.6000 54.8000 144.2000 ;
	    RECT 65.2000 141.6000 66.0000 146.2000 ;
	    RECT 74.8000 141.6000 75.6000 144.2000 ;
	    RECT 78.0000 141.6000 78.8000 144.2000 ;
	    RECT 89.2000 141.6000 90.0000 146.2000 ;
	    RECT 95.6000 141.6000 96.4000 144.2000 ;
	    RECT 100.4000 141.6000 101.2000 146.2000 ;
	    RECT 110.0000 141.6000 110.8000 144.2000 ;
	    RECT 113.2000 141.6000 114.0000 144.2000 ;
	    RECT 124.4000 141.6000 125.2000 146.2000 ;
	    RECT 130.8000 141.6000 131.6000 144.2000 ;
	    RECT 135.6000 141.6000 136.4000 145.4000 ;
	    RECT 140.4000 141.6000 141.2000 144.2000 ;
	    RECT 143.6000 141.6000 144.4000 144.2000 ;
	    RECT 147.8000 141.6000 148.6000 146.0000 ;
	    RECT 153.2000 141.6000 154.0000 146.2000 ;
	    RECT 161.2000 141.6000 162.0000 146.2000 ;
	    RECT 164.4000 141.6000 165.2000 146.2000 ;
	    RECT 167.6000 141.6000 168.4000 146.2000 ;
	    RECT 170.8000 141.6000 171.6000 146.2000 ;
	    RECT 174.0000 141.6000 174.8000 146.2000 ;
	    RECT 176.2000 141.6000 177.0000 146.2000 ;
	    RECT 180.4000 141.6000 181.2000 144.2000 ;
	    RECT 183.6000 141.6000 184.4000 144.2000 ;
	    RECT 188.4000 141.6000 189.2000 146.2000 ;
	    RECT 198.0000 141.6000 198.8000 144.2000 ;
	    RECT 201.2000 141.6000 202.0000 144.2000 ;
	    RECT 212.4000 141.6000 213.2000 146.2000 ;
	    RECT 218.8000 141.6000 219.6000 144.2000 ;
	    RECT 222.0000 141.6000 222.8000 146.2000 ;
	    RECT 0.4000 140.4000 226.8000 141.6000 ;
	    RECT 2.8000 135.8000 3.6000 140.4000 ;
	    RECT 6.0000 137.8000 6.8000 140.4000 ;
	    RECT 10.4000 135.0000 11.2000 140.4000 ;
	    RECT 15.6000 135.4000 16.4000 140.4000 ;
	    RECT 18.8000 137.8000 19.6000 140.4000 ;
	    RECT 25.2000 135.8000 26.0000 140.4000 ;
	    RECT 36.4000 137.8000 37.2000 140.4000 ;
	    RECT 39.6000 137.8000 40.4000 140.4000 ;
	    RECT 49.2000 135.8000 50.0000 140.4000 ;
	    RECT 55.6000 136.6000 56.4000 140.4000 ;
	    RECT 62.0000 135.8000 62.8000 140.4000 ;
	    RECT 71.6000 135.8000 72.4000 140.4000 ;
	    RECT 74.8000 137.8000 75.6000 140.4000 ;
	    RECT 79.0000 135.8000 79.8000 140.4000 ;
	    RECT 82.8000 135.4000 83.6000 140.4000 ;
	    RECT 88.0000 135.0000 88.8000 140.4000 ;
	    RECT 92.4000 137.8000 93.2000 140.4000 ;
	    RECT 94.0000 135.8000 94.8000 140.4000 ;
	    RECT 97.2000 135.8000 98.0000 140.4000 ;
	    RECT 100.4000 135.8000 101.2000 140.4000 ;
	    RECT 103.6000 135.8000 104.4000 140.4000 ;
	    RECT 106.8000 135.8000 107.6000 140.4000 ;
	    RECT 111.6000 135.8000 112.4000 140.4000 ;
	    RECT 121.2000 137.8000 122.0000 140.4000 ;
	    RECT 124.4000 137.8000 125.2000 140.4000 ;
	    RECT 135.6000 135.8000 136.4000 140.4000 ;
	    RECT 142.0000 137.8000 142.8000 140.4000 ;
	    RECT 143.6000 137.8000 144.4000 140.4000 ;
	    RECT 154.8000 135.8000 155.6000 140.4000 ;
	    RECT 164.4000 137.8000 165.2000 140.4000 ;
	    RECT 167.6000 137.8000 168.4000 140.4000 ;
	    RECT 178.8000 135.8000 179.6000 140.4000 ;
	    RECT 185.2000 137.8000 186.0000 140.4000 ;
	    RECT 190.0000 135.8000 190.8000 140.4000 ;
	    RECT 199.6000 137.8000 200.4000 140.4000 ;
	    RECT 202.8000 137.8000 203.6000 140.4000 ;
	    RECT 214.0000 135.8000 214.8000 140.4000 ;
	    RECT 220.4000 137.8000 221.2000 140.4000 ;
	    RECT 2.8000 101.6000 3.6000 106.2000 ;
	    RECT 7.6000 101.6000 8.4000 106.2000 ;
	    RECT 10.8000 101.6000 11.6000 104.2000 ;
	    RECT 14.0000 101.6000 14.8000 104.2000 ;
	    RECT 17.8000 101.6000 18.6000 106.2000 ;
	    RECT 22.0000 101.6000 22.8000 104.2000 ;
	    RECT 25.2000 101.6000 26.0000 105.4000 ;
	    RECT 30.6000 101.6000 31.4000 106.2000 ;
	    RECT 34.8000 101.6000 35.6000 104.2000 ;
	    RECT 36.4000 101.6000 37.2000 104.2000 ;
	    RECT 42.8000 101.6000 43.6000 106.2000 ;
	    RECT 54.0000 101.6000 54.8000 104.2000 ;
	    RECT 57.2000 101.6000 58.0000 104.2000 ;
	    RECT 66.8000 101.6000 67.6000 106.2000 ;
	    RECT 76.4000 101.6000 77.2000 104.2000 ;
	    RECT 79.6000 101.6000 80.4000 106.2000 ;
	    RECT 82.8000 101.6000 83.6000 106.2000 ;
	    RECT 86.0000 101.6000 86.8000 106.2000 ;
	    RECT 89.2000 101.6000 90.0000 106.2000 ;
	    RECT 92.4000 101.6000 93.2000 106.2000 ;
	    RECT 97.2000 101.6000 98.0000 106.2000 ;
	    RECT 106.8000 101.6000 107.6000 104.2000 ;
	    RECT 110.0000 101.6000 110.8000 104.2000 ;
	    RECT 121.2000 101.6000 122.0000 106.2000 ;
	    RECT 127.6000 101.6000 128.4000 104.2000 ;
	    RECT 129.2000 101.6000 130.0000 108.2000 ;
	    RECT 135.6000 101.6000 136.4000 104.2000 ;
	    RECT 138.8000 101.6000 139.6000 104.2000 ;
	    RECT 142.0000 101.6000 142.8000 104.2000 ;
	    RECT 145.2000 101.6000 146.0000 104.2000 ;
	    RECT 150.0000 101.6000 150.8000 105.4000 ;
	    RECT 153.2000 101.6000 154.0000 104.2000 ;
	    RECT 156.4000 101.6000 157.2000 104.2000 ;
	    RECT 163.4000 101.6000 164.2000 106.2000 ;
	    RECT 167.6000 101.6000 168.4000 104.2000 ;
	    RECT 170.8000 101.6000 171.6000 105.4000 ;
	    RECT 175.6000 101.6000 176.4000 106.2000 ;
	    RECT 181.6000 101.6000 182.4000 106.2000 ;
	    RECT 185.2000 101.6000 186.0000 104.2000 ;
	    RECT 188.4000 101.6000 189.2000 106.2000 ;
	    RECT 194.8000 101.6000 195.6000 105.4000 ;
	    RECT 201.2000 101.6000 202.0000 105.4000 ;
	    RECT 204.4000 101.6000 205.2000 106.2000 ;
	    RECT 209.8000 101.6000 210.6000 106.2000 ;
	    RECT 214.0000 101.6000 214.8000 104.2000 ;
	    RECT 217.2000 101.6000 218.0000 104.2000 ;
	    RECT 220.4000 101.6000 221.2000 106.2000 ;
	    RECT 0.4000 100.4000 226.8000 101.6000 ;
	    RECT 1.2000 97.8000 2.0000 100.4000 ;
	    RECT 7.6000 95.8000 8.4000 100.4000 ;
	    RECT 18.8000 97.8000 19.6000 100.4000 ;
	    RECT 22.0000 97.8000 22.8000 100.4000 ;
	    RECT 31.6000 95.8000 32.4000 100.4000 ;
	    RECT 38.0000 95.8000 38.8000 100.4000 ;
	    RECT 44.4000 96.6000 45.2000 100.4000 ;
	    RECT 49.2000 96.4000 50.2000 100.4000 ;
	    RECT 55.4000 99.8000 56.2000 100.4000 ;
	    RECT 55.4000 96.4000 56.4000 99.8000 ;
	    RECT 60.4000 95.8000 61.2000 100.4000 ;
	    RECT 68.4000 97.8000 69.2000 100.4000 ;
	    RECT 74.8000 95.8000 75.6000 100.4000 ;
	    RECT 86.0000 97.8000 86.8000 100.4000 ;
	    RECT 89.2000 97.8000 90.0000 100.4000 ;
	    RECT 98.8000 95.8000 99.6000 100.4000 ;
	    RECT 105.2000 95.8000 106.0000 100.4000 ;
	    RECT 110.0000 95.8000 110.8000 100.4000 ;
	    RECT 114.8000 95.8000 115.6000 100.4000 ;
	    RECT 122.8000 93.8000 123.6000 100.4000 ;
	    RECT 124.4000 93.8000 125.2000 100.4000 ;
	    RECT 132.4000 97.8000 133.2000 100.4000 ;
	    RECT 134.0000 97.8000 134.8000 100.4000 ;
	    RECT 140.4000 95.8000 141.2000 100.4000 ;
	    RECT 151.6000 97.8000 152.4000 100.4000 ;
	    RECT 154.8000 97.8000 155.6000 100.4000 ;
	    RECT 164.4000 95.8000 165.2000 100.4000 ;
	    RECT 177.2000 95.8000 178.0000 100.4000 ;
	    RECT 186.8000 97.8000 187.6000 100.4000 ;
	    RECT 190.0000 97.8000 190.8000 100.4000 ;
	    RECT 201.2000 95.8000 202.0000 100.4000 ;
	    RECT 207.6000 97.8000 208.4000 100.4000 ;
	    RECT 212.4000 95.8000 213.2000 100.4000 ;
	    RECT 215.6000 96.6000 216.4000 100.4000 ;
	    RECT 220.4000 93.8000 221.2000 100.4000 ;
	    RECT 1.2000 61.6000 2.0000 64.2000 ;
	    RECT 7.6000 61.6000 8.4000 66.2000 ;
	    RECT 18.8000 61.6000 19.6000 64.2000 ;
	    RECT 22.0000 61.6000 22.8000 64.2000 ;
	    RECT 31.6000 61.6000 32.4000 66.2000 ;
	    RECT 38.0000 61.6000 38.8000 65.4000 ;
	    RECT 46.0000 61.6000 46.8000 65.4000 ;
	    RECT 49.8000 61.6000 50.6000 66.2000 ;
	    RECT 54.0000 61.6000 54.8000 64.2000 ;
	    RECT 57.2000 61.6000 58.0000 65.4000 ;
	    RECT 66.8000 61.6000 67.6000 64.2000 ;
	    RECT 70.0000 61.6000 70.8000 64.2000 ;
	    RECT 73.2000 61.6000 74.0000 64.2000 ;
	    RECT 78.0000 61.6000 78.8000 65.4000 ;
	    RECT 84.4000 61.6000 85.2000 66.2000 ;
	    RECT 94.0000 61.6000 94.8000 64.2000 ;
	    RECT 97.2000 61.6000 98.0000 64.2000 ;
	    RECT 108.4000 61.6000 109.2000 66.2000 ;
	    RECT 114.8000 61.6000 115.6000 64.2000 ;
	    RECT 116.4000 61.6000 117.2000 64.2000 ;
	    RECT 121.2000 61.6000 122.0000 64.2000 ;
	    RECT 123.2000 61.6000 124.0000 66.2000 ;
	    RECT 129.2000 61.6000 130.0000 66.2000 ;
	    RECT 132.4000 61.6000 133.2000 64.2000 ;
	    RECT 135.6000 61.6000 136.4000 63.8000 ;
	    RECT 151.6000 61.6000 152.4000 66.2000 ;
	    RECT 161.2000 61.6000 162.0000 64.2000 ;
	    RECT 164.4000 61.6000 165.2000 64.2000 ;
	    RECT 175.6000 61.6000 176.4000 66.2000 ;
	    RECT 182.0000 61.6000 182.8000 64.2000 ;
	    RECT 185.2000 61.6000 186.0000 65.4000 ;
	    RECT 191.6000 61.6000 192.4000 65.4000 ;
	    RECT 196.4000 61.6000 197.2000 64.2000 ;
	    RECT 200.6000 61.6000 201.4000 66.2000 ;
	    RECT 206.0000 61.6000 206.8000 65.4000 ;
	    RECT 209.2000 61.6000 210.0000 68.2000 ;
	    RECT 217.2000 61.6000 218.0000 65.4000 ;
	    RECT 222.0000 61.6000 222.8000 64.2000 ;
	    RECT 225.2000 61.6000 226.0000 64.2000 ;
	    RECT 0.4000 60.4000 226.8000 61.6000 ;
	    RECT 2.8000 55.8000 3.6000 60.4000 ;
	    RECT 7.6000 55.8000 8.4000 60.4000 ;
	    RECT 12.0000 55.0000 12.8000 60.4000 ;
	    RECT 17.2000 55.4000 18.0000 60.4000 ;
	    RECT 22.0000 57.8000 22.8000 60.4000 ;
	    RECT 24.2000 55.8000 25.0000 60.4000 ;
	    RECT 28.4000 57.8000 29.2000 60.4000 ;
	    RECT 30.6000 55.8000 31.4000 60.4000 ;
	    RECT 34.8000 57.8000 35.6000 60.4000 ;
	    RECT 38.0000 57.8000 38.8000 60.4000 ;
	    RECT 41.2000 56.4000 42.2000 60.4000 ;
	    RECT 47.4000 59.8000 48.2000 60.4000 ;
	    RECT 47.4000 56.4000 48.4000 59.8000 ;
	    RECT 52.4000 55.4000 53.2000 60.4000 ;
	    RECT 57.6000 55.0000 58.4000 60.4000 ;
	    RECT 62.0000 55.8000 62.8000 60.4000 ;
	    RECT 71.6000 57.8000 72.4000 60.4000 ;
	    RECT 73.2000 55.8000 74.0000 60.4000 ;
	    RECT 76.4000 55.8000 77.2000 60.4000 ;
	    RECT 79.6000 55.8000 80.4000 60.4000 ;
	    RECT 82.8000 55.8000 83.6000 60.4000 ;
	    RECT 86.0000 55.8000 86.8000 60.4000 ;
	    RECT 87.6000 55.8000 88.4000 60.4000 ;
	    RECT 90.8000 55.8000 91.6000 60.4000 ;
	    RECT 94.0000 55.8000 94.8000 60.4000 ;
	    RECT 97.2000 55.8000 98.0000 60.4000 ;
	    RECT 100.4000 55.8000 101.2000 60.4000 ;
	    RECT 102.0000 57.8000 102.8000 60.4000 ;
	    RECT 105.2000 57.8000 106.0000 60.4000 ;
	    RECT 110.0000 55.8000 110.8000 60.4000 ;
	    RECT 111.6000 53.8000 112.4000 60.4000 ;
	    RECT 122.8000 53.8000 123.6000 60.4000 ;
	    RECT 124.4000 57.8000 125.2000 60.4000 ;
	    RECT 130.8000 55.8000 131.6000 60.4000 ;
	    RECT 142.0000 57.8000 142.8000 60.4000 ;
	    RECT 145.2000 57.8000 146.0000 60.4000 ;
	    RECT 154.8000 55.8000 155.6000 60.4000 ;
	    RECT 166.0000 56.6000 166.8000 60.4000 ;
	    RECT 173.4000 56.0000 174.2000 60.4000 ;
	    RECT 180.4000 56.6000 181.2000 60.4000 ;
	    RECT 183.6000 57.8000 184.4000 60.4000 ;
	    RECT 186.8000 57.8000 187.6000 60.4000 ;
	    RECT 190.2000 59.8000 191.0000 60.4000 ;
	    RECT 190.0000 56.4000 191.0000 59.8000 ;
	    RECT 196.2000 56.4000 197.2000 60.4000 ;
	    RECT 202.8000 56.6000 203.6000 60.4000 ;
	    RECT 207.6000 55.8000 208.4000 60.4000 ;
	    RECT 210.8000 57.8000 211.6000 60.4000 ;
	    RECT 214.0000 57.8000 214.8000 60.4000 ;
	    RECT 217.2000 57.8000 218.0000 60.4000 ;
	    RECT 222.0000 55.8000 222.8000 60.4000 ;
	    RECT 1.2000 21.6000 2.0000 24.2000 ;
	    RECT 4.4000 21.6000 5.2000 24.2000 ;
	    RECT 10.8000 21.6000 11.6000 26.2000 ;
	    RECT 22.0000 21.6000 22.8000 24.2000 ;
	    RECT 25.2000 21.6000 26.0000 24.2000 ;
	    RECT 34.8000 21.6000 35.6000 26.2000 ;
	    RECT 42.8000 21.6000 43.6000 26.2000 ;
	    RECT 52.4000 21.6000 53.2000 24.2000 ;
	    RECT 55.6000 21.6000 56.4000 24.2000 ;
	    RECT 66.8000 21.6000 67.6000 26.2000 ;
	    RECT 73.2000 21.6000 74.0000 24.2000 ;
	    RECT 79.6000 21.6000 80.4000 26.2000 ;
	    RECT 87.6000 21.6000 88.4000 25.4000 ;
	    RECT 92.4000 21.6000 93.2000 25.4000 ;
	    RECT 97.2000 21.6000 98.0000 24.2000 ;
	    RECT 100.4000 21.6000 101.2000 28.2000 ;
	    RECT 111.6000 21.6000 112.4000 28.2000 ;
	    RECT 115.4000 21.6000 116.2000 26.0000 ;
	    RECT 119.6000 21.6000 120.4000 24.2000 ;
	    RECT 122.8000 21.6000 123.6000 24.2000 ;
	    RECT 124.4000 21.6000 125.2000 24.2000 ;
	    RECT 130.8000 21.6000 131.6000 26.2000 ;
	    RECT 142.0000 21.6000 142.8000 24.2000 ;
	    RECT 145.2000 21.6000 146.0000 24.2000 ;
	    RECT 154.8000 21.6000 155.6000 26.2000 ;
	    RECT 164.4000 21.6000 165.2000 24.2000 ;
	    RECT 167.6000 21.6000 168.4000 26.2000 ;
	    RECT 172.4000 21.6000 173.2000 24.2000 ;
	    RECT 175.6000 21.6000 176.4000 24.2000 ;
	    RECT 177.2000 21.6000 178.0000 24.2000 ;
	    RECT 182.0000 21.6000 182.8000 25.4000 ;
	    RECT 190.0000 21.6000 190.8000 26.2000 ;
	    RECT 191.6000 21.6000 192.4000 28.2000 ;
	    RECT 201.2000 21.6000 202.0000 25.4000 ;
	    RECT 204.4000 21.6000 205.2000 24.2000 ;
	    RECT 210.8000 21.6000 211.6000 25.4000 ;
	    RECT 214.0000 21.6000 214.8000 28.2000 ;
	    RECT 220.4000 21.6000 221.2000 24.2000 ;
	    RECT 223.6000 21.6000 224.4000 24.2000 ;
	    RECT 0.4000 20.4000 226.8000 21.6000 ;
	    RECT 2.8000 15.8000 3.6000 20.4000 ;
	    RECT 6.0000 17.8000 6.8000 20.4000 ;
	    RECT 12.4000 15.8000 13.2000 20.4000 ;
	    RECT 23.6000 17.8000 24.4000 20.4000 ;
	    RECT 26.8000 17.8000 27.6000 20.4000 ;
	    RECT 36.4000 15.8000 37.2000 20.4000 ;
	    RECT 44.4000 15.8000 45.2000 20.4000 ;
	    RECT 54.0000 17.8000 54.8000 20.4000 ;
	    RECT 57.2000 17.8000 58.0000 20.4000 ;
	    RECT 68.4000 15.8000 69.2000 20.4000 ;
	    RECT 74.8000 17.8000 75.6000 20.4000 ;
	    RECT 82.8000 15.8000 83.6000 20.4000 ;
	    RECT 87.6000 15.8000 88.4000 20.4000 ;
	    RECT 90.8000 17.8000 91.6000 20.4000 ;
	    RECT 97.2000 15.8000 98.0000 20.4000 ;
	    RECT 108.4000 17.8000 109.2000 20.4000 ;
	    RECT 111.6000 17.8000 112.4000 20.4000 ;
	    RECT 121.2000 15.8000 122.0000 20.4000 ;
	    RECT 127.6000 15.8000 128.4000 20.4000 ;
	    RECT 132.4000 15.8000 133.2000 20.4000 ;
	    RECT 135.6000 17.8000 136.4000 20.4000 ;
	    RECT 138.8000 17.8000 139.6000 20.4000 ;
	    RECT 143.0000 16.0000 143.8000 20.4000 ;
	    RECT 148.4000 16.6000 149.2000 20.4000 ;
	    RECT 156.4000 16.6000 157.2000 20.4000 ;
	    RECT 166.0000 15.8000 166.8000 20.4000 ;
	    RECT 169.2000 17.8000 170.0000 20.4000 ;
	    RECT 175.6000 15.8000 176.4000 20.4000 ;
	    RECT 186.8000 17.8000 187.6000 20.4000 ;
	    RECT 190.0000 17.8000 190.8000 20.4000 ;
	    RECT 199.6000 15.8000 200.4000 20.4000 ;
	    RECT 206.0000 16.6000 206.8000 20.4000 ;
	    RECT 212.4000 17.8000 213.2000 20.4000 ;
	    RECT 215.6000 17.8000 216.4000 20.4000 ;
	    RECT 218.8000 17.8000 219.6000 20.4000 ;
	    RECT 222.0000 15.8000 222.8000 20.4000 ;
         LAYER metal2 ;
	    RECT 154.4000 180.6000 159.2000 181.4000 ;
	    RECT 154.4000 140.6000 159.2000 141.4000 ;
	    RECT 154.4000 100.6000 159.2000 101.4000 ;
	    RECT 154.4000 60.6000 159.2000 61.4000 ;
	    RECT 154.4000 20.6000 159.2000 21.4000 ;
         LAYER metal3 ;
	    RECT 154.4000 180.4000 159.2000 181.6000 ;
	    RECT 154.4000 140.4000 159.2000 141.6000 ;
	    RECT 154.4000 100.4000 159.2000 101.6000 ;
	    RECT 154.4000 60.4000 159.2000 61.6000 ;
	    RECT 154.4000 20.4000 159.2000 21.6000 ;
         LAYER metal4 ;
	    RECT 154.4000 -4.0000 159.2000 204.0000 ;
      END
   END gnd
   PIN clock
      PORT
         LAYER metal1 ;
	    RECT 161.2000 148.2000 163.0000 149.0000 ;
	    RECT 161.2000 147.6000 162.0000 148.2000 ;
	    RECT 106.8000 133.8000 107.6000 134.4000 ;
	    RECT 105.8000 133.0000 107.6000 133.8000 ;
	    RECT 91.4000 108.2000 93.2000 109.0000 ;
	    RECT 92.4000 107.6000 93.2000 108.2000 ;
	    RECT 86.0000 54.3000 86.8000 54.4000 ;
	    RECT 87.6000 54.3000 88.4000 54.4000 ;
	    RECT 86.0000 53.8000 88.4000 54.3000 ;
	    RECT 85.0000 53.7000 89.4000 53.8000 ;
	    RECT 85.0000 53.0000 86.8000 53.7000 ;
	    RECT 87.6000 53.0000 89.4000 53.7000 ;
         LAYER metal2 ;
	    RECT 161.2000 148.3000 162.0000 148.4000 ;
	    RECT 162.9000 148.3000 163.5000 204.3000 ;
	    RECT 161.2000 147.7000 163.5000 148.3000 ;
	    RECT 161.2000 147.6000 162.0000 147.7000 ;
	    RECT 106.8000 133.6000 107.6000 134.4000 ;
	    RECT 106.9000 130.4000 107.5000 133.6000 ;
	    RECT 92.4000 129.6000 93.2000 130.4000 ;
	    RECT 106.8000 129.6000 107.6000 130.4000 ;
	    RECT 92.5000 108.4000 93.1000 129.6000 ;
	    RECT 92.4000 107.6000 93.2000 108.4000 ;
	    RECT 92.5000 100.4000 93.1000 107.6000 ;
	    RECT 92.4000 99.6000 93.2000 100.4000 ;
	    RECT 87.6000 59.6000 88.4000 60.4000 ;
	    RECT 87.7000 54.4000 88.3000 59.6000 ;
	    RECT 87.6000 53.6000 88.4000 54.4000 ;
         LAYER metal3 ;
	    RECT 151.6000 148.3000 152.4000 148.4000 ;
	    RECT 161.2000 148.3000 162.0000 148.4000 ;
	    RECT 151.6000 147.7000 162.0000 148.3000 ;
	    RECT 151.6000 147.6000 152.4000 147.7000 ;
	    RECT 161.2000 147.6000 162.0000 147.7000 ;
	    RECT 92.4000 130.3000 93.2000 130.4000 ;
	    RECT 106.8000 130.3000 107.6000 130.4000 ;
	    RECT 151.6000 130.3000 152.4000 130.4000 ;
	    RECT 92.4000 129.7000 152.4000 130.3000 ;
	    RECT 92.4000 129.6000 93.2000 129.7000 ;
	    RECT 106.8000 129.6000 107.6000 129.7000 ;
	    RECT 151.6000 129.6000 152.4000 129.7000 ;
	    RECT 87.6000 100.3000 88.4000 100.4000 ;
	    RECT 92.4000 100.3000 93.2000 100.4000 ;
	    RECT 87.6000 99.7000 93.2000 100.3000 ;
	    RECT 87.6000 99.6000 88.4000 99.7000 ;
	    RECT 92.4000 99.6000 93.2000 99.7000 ;
	    RECT 87.6000 59.6000 88.4000 60.4000 ;
         LAYER metal4 ;
	    RECT 151.4000 129.4000 152.6000 148.6000 ;
	    RECT 87.4000 59.4000 88.6000 100.6000 ;
      END
   END clock
   PIN reset
      PORT
         LAYER metal1 ;
	    RECT 138.8000 175.6000 139.6000 177.2000 ;
         LAYER metal2 ;
	    RECT 137.3000 203.7000 139.5000 204.3000 ;
	    RECT 138.9000 176.4000 139.5000 203.7000 ;
	    RECT 138.8000 175.6000 139.6000 176.4000 ;
      END
   END reset
   PIN start
      PORT
         LAYER metal1 ;
	    RECT 186.8000 186.8000 187.6000 188.4000 ;
         LAYER metal2 ;
	    RECT 182.1000 200.4000 182.7000 204.3000 ;
	    RECT 182.0000 199.6000 182.8000 200.4000 ;
	    RECT 186.8000 199.6000 187.6000 200.4000 ;
	    RECT 186.9000 188.4000 187.5000 199.6000 ;
	    RECT 186.8000 187.6000 187.6000 188.4000 ;
         LAYER metal3 ;
	    RECT 182.0000 200.3000 182.8000 200.4000 ;
	    RECT 186.8000 200.3000 187.6000 200.4000 ;
	    RECT 182.0000 199.7000 187.6000 200.3000 ;
	    RECT 182.0000 199.6000 182.8000 199.7000 ;
	    RECT 186.8000 199.6000 187.6000 199.7000 ;
      END
   END start
   PIN N[0]
      PORT
         LAYER metal1 ;
	    RECT 201.2000 184.8000 202.0000 186.4000 ;
         LAYER metal2 ;
	    RECT 201.3000 203.7000 203.5000 204.3000 ;
	    RECT 201.3000 186.4000 201.9000 203.7000 ;
	    RECT 201.2000 185.6000 202.0000 186.4000 ;
      END
   END N[0]
   PIN N[1]
      PORT
         LAYER metal1 ;
	    RECT 214.0000 55.6000 214.8000 57.2000 ;
	    RECT 222.0000 53.6000 222.8000 55.2000 ;
	    RECT 212.4000 15.6000 213.2000 17.2000 ;
         LAYER metal2 ;
	    RECT 214.0000 57.6000 214.8000 58.4000 ;
	    RECT 222.0000 57.6000 222.8000 58.4000 ;
	    RECT 214.1000 56.4000 214.7000 57.6000 ;
	    RECT 214.0000 56.3000 214.8000 56.4000 ;
	    RECT 212.5000 55.7000 214.8000 56.3000 ;
	    RECT 212.5000 16.4000 213.1000 55.7000 ;
	    RECT 214.0000 55.6000 214.8000 55.7000 ;
	    RECT 222.1000 54.4000 222.7000 57.6000 ;
	    RECT 222.0000 53.6000 222.8000 54.4000 ;
	    RECT 212.4000 15.6000 213.2000 16.4000 ;
         LAYER metal3 ;
	    RECT 214.0000 58.3000 214.8000 58.4000 ;
	    RECT 222.0000 58.3000 222.8000 58.4000 ;
	    RECT 214.0000 57.7000 229.1000 58.3000 ;
	    RECT 214.0000 57.6000 214.8000 57.7000 ;
	    RECT 222.0000 57.6000 222.8000 57.7000 ;
      END
   END N[1]
   PIN N[2]
      PORT
         LAYER metal1 ;
	    RECT 217.2000 52.3000 218.0000 52.4000 ;
	    RECT 218.8000 52.3000 219.6000 52.4000 ;
	    RECT 217.2000 51.7000 219.6000 52.3000 ;
	    RECT 217.2000 50.8000 218.0000 51.7000 ;
	    RECT 218.8000 51.6000 219.6000 51.7000 ;
	    RECT 218.9000 50.4000 219.5000 51.6000 ;
	    RECT 218.8000 48.8000 219.6000 50.4000 ;
         LAYER metal2 ;
	    RECT 218.8000 53.6000 219.6000 54.4000 ;
	    RECT 218.9000 52.4000 219.5000 53.6000 ;
	    RECT 218.8000 51.6000 219.6000 52.4000 ;
         LAYER metal3 ;
	    RECT 218.8000 54.3000 219.6000 54.4000 ;
	    RECT 218.8000 53.7000 229.1000 54.3000 ;
	    RECT 218.8000 53.6000 219.6000 53.7000 ;
      END
   END N[2]
   PIN N[3]
      PORT
         LAYER metal1 ;
	    RECT 199.6000 67.6000 200.4000 69.2000 ;
	    RECT 207.6000 68.2000 208.4000 68.4000 ;
	    RECT 206.8000 67.6000 208.4000 68.2000 ;
	    RECT 215.6000 68.2000 216.4000 68.4000 ;
	    RECT 215.6000 67.6000 217.2000 68.2000 ;
	    RECT 206.8000 67.2000 207.6000 67.6000 ;
	    RECT 216.4000 67.2000 217.2000 67.6000 ;
	    RECT 225.2000 64.8000 226.0000 66.4000 ;
         LAYER metal2 ;
	    RECT 199.6000 67.6000 200.4000 68.4000 ;
	    RECT 207.6000 67.6000 208.4000 68.4000 ;
	    RECT 215.6000 67.6000 216.4000 68.4000 ;
	    RECT 225.2000 67.6000 226.0000 68.4000 ;
	    RECT 225.3000 66.4000 225.9000 67.6000 ;
	    RECT 225.2000 65.6000 226.0000 66.4000 ;
         LAYER metal3 ;
	    RECT 199.6000 68.3000 200.4000 68.4000 ;
	    RECT 207.6000 68.3000 208.4000 68.4000 ;
	    RECT 215.6000 68.3000 216.4000 68.4000 ;
	    RECT 225.2000 68.3000 226.0000 68.4000 ;
	    RECT 199.6000 67.7000 229.1000 68.3000 ;
	    RECT 199.6000 67.6000 200.4000 67.7000 ;
	    RECT 207.6000 67.6000 208.4000 67.7000 ;
	    RECT 215.6000 67.6000 216.4000 67.7000 ;
	    RECT 225.2000 67.6000 226.0000 67.7000 ;
      END
   END N[3]
   PIN N[4]
      PORT
         LAYER metal1 ;
	    RECT 219.6000 73.6000 220.4000 74.4000 ;
	    RECT 219.8000 72.4000 220.4000 73.6000 ;
	    RECT 219.8000 71.8000 221.2000 72.4000 ;
	    RECT 220.4000 71.6000 221.2000 71.8000 ;
	    RECT 220.5000 70.3000 221.1000 71.6000 ;
	    RECT 222.0000 70.3000 222.8000 71.2000 ;
	    RECT 220.5000 69.7000 222.8000 70.3000 ;
	    RECT 222.0000 69.6000 222.8000 69.7000 ;
         LAYER metal2 ;
	    RECT 220.4000 71.6000 221.2000 72.4000 ;
         LAYER metal3 ;
	    RECT 220.4000 72.3000 221.2000 72.4000 ;
	    RECT 220.4000 71.7000 229.1000 72.3000 ;
	    RECT 220.4000 71.6000 221.2000 71.7000 ;
      END
   END N[4]
   PIN N[5]
      PORT
         LAYER metal1 ;
	    RECT 202.8000 108.2000 203.6000 108.4000 ;
	    RECT 202.0000 107.6000 203.6000 108.2000 ;
	    RECT 202.0000 107.2000 202.8000 107.6000 ;
	    RECT 217.2000 104.8000 218.0000 106.4000 ;
	    RECT 214.8000 94.4000 215.6000 94.8000 ;
	    RECT 214.0000 93.8000 215.6000 94.4000 ;
	    RECT 214.0000 93.6000 214.8000 93.8000 ;
	    RECT 220.4000 24.8000 221.2000 26.4000 ;
         LAYER metal2 ;
	    RECT 202.8000 107.6000 203.6000 108.4000 ;
	    RECT 202.9000 96.4000 203.5000 107.6000 ;
	    RECT 217.2000 105.6000 218.0000 106.4000 ;
	    RECT 217.3000 96.4000 217.9000 105.6000 ;
	    RECT 202.8000 95.6000 203.6000 96.4000 ;
	    RECT 214.0000 95.6000 214.8000 96.4000 ;
	    RECT 217.2000 95.6000 218.0000 96.4000 ;
	    RECT 214.1000 94.4000 214.7000 95.6000 ;
	    RECT 214.0000 93.6000 214.8000 94.4000 ;
	    RECT 220.4000 25.6000 221.2000 26.4000 ;
         LAYER metal3 ;
	    RECT 202.8000 96.3000 203.6000 96.4000 ;
	    RECT 214.0000 96.3000 214.8000 96.4000 ;
	    RECT 217.2000 96.3000 218.0000 96.4000 ;
	    RECT 225.2000 96.3000 226.0000 96.4000 ;
	    RECT 202.8000 95.7000 226.0000 96.3000 ;
	    RECT 202.8000 95.6000 203.6000 95.7000 ;
	    RECT 214.0000 95.6000 214.8000 95.7000 ;
	    RECT 217.2000 95.6000 218.0000 95.7000 ;
	    RECT 225.2000 95.6000 226.0000 95.7000 ;
	    RECT 220.4000 26.3000 221.2000 26.4000 ;
	    RECT 225.2000 26.3000 226.0000 26.4000 ;
	    RECT 220.4000 25.7000 229.1000 26.3000 ;
	    RECT 220.4000 25.6000 221.2000 25.7000 ;
	    RECT 225.2000 25.6000 226.0000 25.7000 ;
         LAYER metal4 ;
	    RECT 225.0000 25.4000 226.2000 96.6000 ;
      END
   END N[5]
   PIN N[6]
      PORT
         LAYER metal1 ;
	    RECT 218.8000 90.2000 219.6000 90.4000 ;
	    RECT 218.2000 89.6000 219.6000 90.2000 ;
	    RECT 218.2000 88.4000 218.8000 89.6000 ;
	    RECT 218.0000 88.3000 218.8000 88.4000 ;
	    RECT 220.4000 88.3000 221.2000 88.4000 ;
	    RECT 218.0000 87.7000 221.2000 88.3000 ;
	    RECT 218.0000 87.6000 218.8000 87.7000 ;
	    RECT 220.4000 87.6000 221.2000 87.7000 ;
	    RECT 223.6000 30.3000 224.4000 31.2000 ;
	    RECT 225.2000 30.3000 226.0000 30.4000 ;
	    RECT 223.6000 29.7000 226.0000 30.3000 ;
	    RECT 223.6000 29.6000 224.4000 29.7000 ;
	    RECT 225.2000 29.6000 226.0000 29.7000 ;
         LAYER metal2 ;
	    RECT 220.4000 87.6000 221.2000 88.4000 ;
	    RECT 220.5000 86.4000 221.1000 87.6000 ;
	    RECT 220.4000 85.6000 221.2000 86.4000 ;
	    RECT 225.2000 33.6000 226.0000 34.4000 ;
	    RECT 225.3000 30.4000 225.9000 33.6000 ;
	    RECT 225.2000 29.6000 226.0000 30.4000 ;
         LAYER metal3 ;
	    RECT 220.4000 86.3000 221.2000 86.4000 ;
	    RECT 222.0000 86.3000 222.8000 86.4000 ;
	    RECT 220.4000 85.7000 222.8000 86.3000 ;
	    RECT 220.4000 85.6000 221.2000 85.7000 ;
	    RECT 222.0000 85.6000 222.8000 85.7000 ;
	    RECT 222.0000 34.3000 222.8000 34.4000 ;
	    RECT 225.2000 34.3000 226.0000 34.4000 ;
	    RECT 222.0000 33.7000 229.1000 34.3000 ;
	    RECT 222.0000 33.6000 222.8000 33.7000 ;
	    RECT 225.2000 33.6000 226.0000 33.7000 ;
         LAYER metal4 ;
	    RECT 221.8000 33.4000 223.0000 86.6000 ;
      END
   END N[6]
   PIN N[7]
      PORT
         LAYER metal1 ;
	    RECT 222.0000 186.3000 222.8000 186.4000 ;
	    RECT 225.2000 186.3000 226.0000 186.4000 ;
	    RECT 222.0000 185.7000 226.0000 186.3000 ;
	    RECT 222.0000 184.8000 222.8000 185.7000 ;
	    RECT 225.2000 185.6000 226.0000 185.7000 ;
	    RECT 202.8000 28.2000 203.6000 28.4000 ;
	    RECT 202.0000 27.6000 203.6000 28.2000 ;
	    RECT 202.0000 27.2000 202.8000 27.6000 ;
	    RECT 205.2000 14.4000 206.0000 14.8000 ;
	    RECT 204.4000 13.8000 206.0000 14.4000 ;
	    RECT 204.4000 13.6000 205.2000 13.8000 ;
         LAYER metal2 ;
	    RECT 215.6000 185.6000 216.4000 186.4000 ;
	    RECT 225.2000 185.6000 226.0000 186.4000 ;
	    RECT 215.7000 94.4000 216.3000 185.6000 ;
	    RECT 215.6000 93.6000 216.4000 94.4000 ;
	    RECT 202.8000 27.6000 203.6000 28.4000 ;
	    RECT 202.9000 14.3000 203.5000 27.6000 ;
	    RECT 204.4000 14.3000 205.2000 14.4000 ;
	    RECT 202.9000 13.7000 205.2000 14.3000 ;
	    RECT 204.4000 13.6000 205.2000 13.7000 ;
         LAYER metal3 ;
	    RECT 215.6000 186.3000 216.4000 186.4000 ;
	    RECT 225.2000 186.3000 226.0000 186.4000 ;
	    RECT 215.6000 185.7000 229.1000 186.3000 ;
	    RECT 215.6000 185.6000 216.4000 185.7000 ;
	    RECT 225.2000 185.6000 226.0000 185.7000 ;
	    RECT 215.6000 93.6000 216.4000 94.4000 ;
	    RECT 202.8000 28.3000 203.6000 28.4000 ;
	    RECT 215.6000 28.3000 216.4000 28.4000 ;
	    RECT 202.8000 27.7000 216.4000 28.3000 ;
	    RECT 202.8000 27.6000 203.6000 27.7000 ;
	    RECT 215.6000 27.6000 216.4000 27.7000 ;
         LAYER metal4 ;
	    RECT 215.4000 27.4000 216.6000 94.6000 ;
      END
   END N[7]
   PIN N[8]
      PORT
         LAYER metal1 ;
	    RECT 215.6000 29.6000 217.2000 30.4000 ;
	    RECT 215.6000 15.6000 216.4000 17.2000 ;
         LAYER metal2 ;
	    RECT 215.6000 29.6000 216.4000 30.4000 ;
	    RECT 215.7000 26.4000 216.3000 29.6000 ;
	    RECT 215.6000 25.6000 216.4000 26.4000 ;
	    RECT 215.7000 16.4000 216.3000 25.6000 ;
	    RECT 215.6000 15.6000 216.4000 16.4000 ;
         LAYER metal3 ;
	    RECT 218.8000 30.3000 219.6000 30.4000 ;
	    RECT 218.8000 29.7000 229.1000 30.3000 ;
	    RECT 218.8000 29.6000 219.6000 29.7000 ;
	    RECT 215.6000 26.3000 216.4000 26.4000 ;
	    RECT 218.8000 26.3000 219.6000 26.4000 ;
	    RECT 215.6000 25.7000 219.6000 26.3000 ;
	    RECT 215.6000 25.6000 216.4000 25.7000 ;
	    RECT 218.8000 25.6000 219.6000 25.7000 ;
         LAYER metal4 ;
	    RECT 218.6000 25.4000 219.8000 30.6000 ;
      END
   END N[8]
   PIN dp[0]
      PORT
         LAYER metal1 ;
	    RECT 215.6000 191.8000 216.4000 199.8000 ;
	    RECT 215.6000 189.6000 216.2000 191.8000 ;
	    RECT 215.6000 182.2000 216.4000 189.6000 ;
         LAYER metal2 ;
	    RECT 215.7000 203.7000 217.9000 204.3000 ;
	    RECT 215.7000 198.4000 216.3000 203.7000 ;
	    RECT 215.6000 197.6000 216.4000 198.4000 ;
      END
   END dp[0]
   PIN dp[1]
      PORT
         LAYER metal1 ;
	    RECT 86.0000 191.8000 86.8000 199.8000 ;
	    RECT 86.0000 189.6000 86.6000 191.8000 ;
	    RECT 86.0000 182.2000 86.8000 189.6000 ;
         LAYER metal2 ;
	    RECT 86.1000 198.4000 86.7000 204.3000 ;
	    RECT 86.0000 197.6000 86.8000 198.4000 ;
      END
   END dp[1]
   PIN dp[2]
      PORT
         LAYER metal1 ;
	    RECT 41.2000 191.8000 42.0000 199.8000 ;
	    RECT 41.2000 189.6000 41.8000 191.8000 ;
	    RECT 41.2000 182.2000 42.0000 189.6000 ;
         LAYER metal2 ;
	    RECT 41.3000 203.7000 43.5000 204.3000 ;
	    RECT 41.3000 198.4000 41.9000 203.7000 ;
	    RECT 41.2000 197.6000 42.0000 198.4000 ;
      END
   END dp[2]
   PIN dp[3]
      PORT
         LAYER metal1 ;
	    RECT 159.6000 198.3000 160.4000 198.4000 ;
	    RECT 161.2000 198.3000 162.0000 199.8000 ;
	    RECT 159.6000 197.7000 162.0000 198.3000 ;
	    RECT 159.6000 197.6000 160.4000 197.7000 ;
	    RECT 161.2000 191.8000 162.0000 197.7000 ;
	    RECT 161.2000 189.6000 161.8000 191.8000 ;
	    RECT 161.2000 182.2000 162.0000 189.6000 ;
         LAYER metal2 ;
	    RECT 159.7000 198.4000 160.3000 204.3000 ;
	    RECT 159.6000 197.6000 160.4000 198.4000 ;
      END
   END dp[3]
   PIN dp[4]
      PORT
         LAYER metal1 ;
	    RECT 98.8000 191.8000 99.6000 199.8000 ;
	    RECT 99.0000 189.6000 99.6000 191.8000 ;
	    RECT 98.8000 182.2000 99.6000 189.6000 ;
         LAYER metal2 ;
	    RECT 97.3000 203.7000 99.5000 204.3000 ;
	    RECT 98.9000 198.4000 99.5000 203.7000 ;
	    RECT 98.8000 197.6000 99.6000 198.4000 ;
      END
   END dp[4]
   PIN dp[5]
      PORT
         LAYER metal1 ;
	    RECT 1.2000 151.8000 2.0000 159.8000 ;
	    RECT 1.2000 149.6000 1.8000 151.8000 ;
	    RECT 1.2000 142.2000 2.0000 149.6000 ;
         LAYER metal2 ;
	    RECT 1.2000 149.6000 2.0000 150.4000 ;
	    RECT 1.3000 148.4000 1.9000 149.6000 ;
	    RECT 1.2000 147.6000 2.0000 148.4000 ;
         LAYER metal3 ;
	    RECT 1.2000 150.3000 2.0000 150.4000 ;
	    RECT -1.9000 149.7000 2.0000 150.3000 ;
	    RECT 1.2000 149.6000 2.0000 149.7000 ;
      END
   END dp[5]
   PIN dp[6]
      PORT
         LAYER metal1 ;
	    RECT 1.2000 191.8000 2.0000 199.8000 ;
	    RECT 1.2000 189.6000 1.8000 191.8000 ;
	    RECT 1.2000 182.2000 2.0000 189.6000 ;
         LAYER metal2 ;
	    RECT 1.2000 189.6000 2.0000 190.4000 ;
	    RECT 1.3000 188.4000 1.9000 189.6000 ;
	    RECT 1.2000 187.6000 2.0000 188.4000 ;
         LAYER metal3 ;
	    RECT 1.2000 190.3000 2.0000 190.4000 ;
	    RECT -1.9000 189.7000 2.0000 190.3000 ;
	    RECT 1.2000 189.6000 2.0000 189.7000 ;
      END
   END dp[6]
   PIN dp[7]
      PORT
         LAYER metal1 ;
	    RECT 1.2000 12.4000 2.0000 19.8000 ;
	    RECT 1.2000 10.2000 1.8000 12.4000 ;
	    RECT 1.2000 2.2000 2.0000 10.2000 ;
         LAYER metal2 ;
	    RECT 1.2000 9.6000 2.0000 10.4000 ;
	    RECT 1.3000 8.4000 1.9000 9.6000 ;
	    RECT 1.2000 7.6000 2.0000 8.4000 ;
         LAYER metal3 ;
	    RECT 1.2000 10.3000 2.0000 10.4000 ;
	    RECT -1.9000 9.7000 2.0000 10.3000 ;
	    RECT 1.2000 9.6000 2.0000 9.7000 ;
      END
   END dp[7]
   PIN dp[8]
      PORT
         LAYER metal1 ;
	    RECT 84.4000 12.4000 85.2000 19.8000 ;
	    RECT 84.6000 10.2000 85.2000 12.4000 ;
	    RECT 84.4000 2.2000 85.2000 10.2000 ;
         LAYER metal2 ;
	    RECT 84.4000 3.6000 85.2000 4.4000 ;
	    RECT 84.5000 2.4000 85.1000 3.6000 ;
	    RECT 81.2000 1.6000 82.0000 2.4000 ;
	    RECT 84.4000 1.6000 85.2000 2.4000 ;
	    RECT 81.3000 -2.3000 81.9000 1.6000 ;
         LAYER metal3 ;
	    RECT 81.2000 2.3000 82.0000 2.4000 ;
	    RECT 84.4000 2.3000 85.2000 2.4000 ;
	    RECT 81.2000 1.7000 85.2000 2.3000 ;
	    RECT 81.2000 1.6000 82.0000 1.7000 ;
	    RECT 84.4000 1.6000 85.2000 1.7000 ;
      END
   END dp[8]
   PIN done
      PORT
         LAYER metal1 ;
	    RECT 223.6000 151.8000 224.4000 159.8000 ;
	    RECT 223.8000 149.6000 224.4000 151.8000 ;
	    RECT 223.6000 148.3000 224.4000 149.6000 ;
	    RECT 225.2000 148.3000 226.0000 148.4000 ;
	    RECT 223.6000 147.7000 226.0000 148.3000 ;
	    RECT 223.6000 142.2000 224.4000 147.7000 ;
	    RECT 225.2000 147.6000 226.0000 147.7000 ;
         LAYER metal2 ;
	    RECT 225.2000 149.6000 226.0000 150.4000 ;
	    RECT 225.3000 148.4000 225.9000 149.6000 ;
	    RECT 225.2000 147.6000 226.0000 148.4000 ;
         LAYER metal3 ;
	    RECT 225.2000 150.3000 226.0000 150.4000 ;
	    RECT 225.2000 149.7000 229.1000 150.3000 ;
	    RECT 225.2000 149.6000 226.0000 149.7000 ;
      END
   END done
   PIN counter[0]
      PORT
         LAYER metal1 ;
	    RECT 134.0000 12.4000 134.8000 19.8000 ;
	    RECT 134.2000 10.2000 134.8000 12.4000 ;
	    RECT 134.0000 2.2000 134.8000 10.2000 ;
         LAYER metal2 ;
	    RECT 134.0000 3.6000 134.8000 4.4000 ;
	    RECT 134.1000 -1.7000 134.7000 3.6000 ;
	    RECT 132.5000 -2.3000 134.7000 -1.7000 ;
      END
   END counter[0]
   PIN counter[1]
      PORT
         LAYER metal1 ;
	    RECT 164.4000 12.4000 165.2000 19.8000 ;
	    RECT 164.4000 10.2000 165.0000 12.4000 ;
	    RECT 164.4000 2.2000 165.2000 10.2000 ;
         LAYER metal2 ;
	    RECT 164.4000 3.6000 165.2000 4.4000 ;
	    RECT 164.5000 -1.7000 165.1000 3.6000 ;
	    RECT 164.5000 -2.3000 166.7000 -1.7000 ;
      END
   END counter[1]
   PIN counter[2]
      PORT
         LAYER metal1 ;
	    RECT 209.2000 52.4000 210.0000 59.8000 ;
	    RECT 209.4000 50.2000 210.0000 52.4000 ;
	    RECT 209.2000 48.3000 210.0000 50.2000 ;
	    RECT 210.8000 48.3000 211.6000 48.4000 ;
	    RECT 209.2000 47.7000 211.6000 48.3000 ;
	    RECT 209.2000 42.2000 210.0000 47.7000 ;
	    RECT 210.8000 47.6000 211.6000 47.7000 ;
         LAYER metal2 ;
	    RECT 210.8000 49.6000 211.6000 50.4000 ;
	    RECT 210.9000 48.4000 211.5000 49.6000 ;
	    RECT 210.8000 47.6000 211.6000 48.4000 ;
         LAYER metal3 ;
	    RECT 210.8000 50.3000 211.6000 50.4000 ;
	    RECT 210.8000 49.7000 229.1000 50.3000 ;
	    RECT 210.8000 49.6000 211.6000 49.7000 ;
      END
   END counter[2]
   PIN counter[3]
      PORT
         LAYER metal1 ;
	    RECT 223.6000 12.4000 224.4000 19.8000 ;
	    RECT 223.8000 10.2000 224.4000 12.4000 ;
	    RECT 223.6000 8.3000 224.4000 10.2000 ;
	    RECT 225.2000 8.3000 226.0000 8.4000 ;
	    RECT 223.6000 7.7000 226.0000 8.3000 ;
	    RECT 223.6000 2.2000 224.4000 7.7000 ;
	    RECT 225.2000 7.6000 226.0000 7.7000 ;
         LAYER metal2 ;
	    RECT 225.2000 9.6000 226.0000 10.4000 ;
	    RECT 225.3000 8.4000 225.9000 9.6000 ;
	    RECT 225.2000 7.6000 226.0000 8.4000 ;
         LAYER metal3 ;
	    RECT 225.2000 10.3000 226.0000 10.4000 ;
	    RECT 225.2000 9.7000 229.1000 10.3000 ;
	    RECT 225.2000 9.6000 226.0000 9.7000 ;
      END
   END counter[3]
   PIN counter[4]
      PORT
         LAYER metal1 ;
	    RECT 222.0000 114.3000 222.8000 119.8000 ;
	    RECT 225.2000 114.3000 226.0000 114.4000 ;
	    RECT 222.0000 113.7000 226.0000 114.3000 ;
	    RECT 222.0000 111.8000 222.8000 113.7000 ;
	    RECT 225.2000 113.6000 226.0000 113.7000 ;
	    RECT 222.2000 109.6000 222.8000 111.8000 ;
	    RECT 222.0000 102.2000 222.8000 109.6000 ;
         LAYER metal2 ;
	    RECT 225.2000 113.6000 226.0000 114.4000 ;
         LAYER metal3 ;
	    RECT 225.2000 114.3000 226.0000 114.4000 ;
	    RECT 225.2000 113.7000 229.1000 114.3000 ;
	    RECT 225.2000 113.6000 226.0000 113.7000 ;
      END
   END counter[4]
   PIN counter[5]
      PORT
         LAYER metal1 ;
	    RECT 190.0000 111.8000 190.8000 119.8000 ;
	    RECT 190.2000 109.6000 190.8000 111.8000 ;
	    RECT 190.0000 102.2000 190.8000 109.6000 ;
         LAYER metal2 ;
	    RECT 190.0000 113.6000 190.8000 114.4000 ;
	    RECT 190.1000 112.4000 190.7000 113.6000 ;
	    RECT 190.0000 111.6000 190.8000 112.4000 ;
         LAYER metal3 ;
	    RECT 190.0000 112.3000 190.8000 112.4000 ;
	    RECT 190.0000 111.7000 229.1000 112.3000 ;
	    RECT 190.0000 111.6000 190.8000 111.7000 ;
	    RECT 228.5000 109.7000 229.1000 111.7000 ;
      END
   END counter[5]
   PIN counter[6]
      PORT
         LAYER metal1 ;
	    RECT 129.2000 12.4000 130.0000 19.8000 ;
	    RECT 129.4000 10.2000 130.0000 12.4000 ;
	    RECT 129.2000 2.2000 130.0000 10.2000 ;
         LAYER metal2 ;
	    RECT 129.2000 3.6000 130.0000 4.4000 ;
	    RECT 129.3000 -1.7000 129.9000 3.6000 ;
	    RECT 127.7000 -2.3000 129.9000 -1.7000 ;
      END
   END counter[6]
   PIN counter[7]
      PORT
         LAYER metal1 ;
	    RECT 86.0000 12.4000 86.8000 19.8000 ;
	    RECT 86.0000 10.2000 86.6000 12.4000 ;
	    RECT 86.0000 2.2000 86.8000 10.2000 ;
         LAYER metal2 ;
	    RECT 86.0000 3.6000 86.8000 4.4000 ;
	    RECT 86.1000 -1.7000 86.7000 3.6000 ;
	    RECT 86.1000 -2.3000 88.3000 -1.7000 ;
      END
   END counter[7]
   PIN sr[0]
      PORT
         LAYER metal1 ;
	    RECT 94.0000 191.8000 94.8000 199.8000 ;
	    RECT 94.2000 189.6000 94.8000 191.8000 ;
	    RECT 94.0000 182.2000 94.8000 189.6000 ;
         LAYER metal2 ;
	    RECT 92.5000 203.7000 94.7000 204.3000 ;
	    RECT 94.1000 198.4000 94.7000 203.7000 ;
	    RECT 94.0000 197.6000 94.8000 198.4000 ;
      END
   END sr[0]
   PIN sr[1]
      PORT
         LAYER metal1 ;
	    RECT 1.2000 172.4000 2.0000 179.8000 ;
	    RECT 1.2000 170.2000 1.8000 172.4000 ;
	    RECT 1.2000 162.2000 2.0000 170.2000 ;
         LAYER metal2 ;
	    RECT 1.2000 169.6000 2.0000 170.4000 ;
	    RECT 1.3000 168.4000 1.9000 169.6000 ;
	    RECT 1.2000 167.6000 2.0000 168.4000 ;
         LAYER metal3 ;
	    RECT 1.2000 170.3000 2.0000 170.4000 ;
	    RECT -1.9000 169.7000 2.0000 170.3000 ;
	    RECT 1.2000 169.6000 2.0000 169.7000 ;
      END
   END sr[1]
   PIN sr[2]
      PORT
         LAYER metal1 ;
	    RECT 1.2000 132.4000 2.0000 139.8000 ;
	    RECT 1.2000 130.2000 1.8000 132.4000 ;
	    RECT 1.2000 122.2000 2.0000 130.2000 ;
         LAYER metal2 ;
	    RECT 1.2000 129.6000 2.0000 130.4000 ;
	    RECT 1.3000 128.4000 1.9000 129.6000 ;
	    RECT 1.2000 127.6000 2.0000 128.4000 ;
         LAYER metal3 ;
	    RECT 1.2000 130.3000 2.0000 130.4000 ;
	    RECT -1.9000 129.7000 2.0000 130.3000 ;
	    RECT 1.2000 129.6000 2.0000 129.7000 ;
      END
   END sr[2]
   PIN sr[3]
      PORT
         LAYER metal1 ;
	    RECT 36.4000 92.4000 37.2000 99.8000 ;
	    RECT 36.4000 90.2000 37.0000 92.4000 ;
	    RECT 36.4000 82.2000 37.2000 90.2000 ;
         LAYER metal2 ;
	    RECT 36.4000 93.6000 37.2000 94.4000 ;
	    RECT 36.5000 90.4000 37.1000 93.6000 ;
	    RECT 36.4000 89.6000 37.2000 90.4000 ;
         LAYER metal3 ;
	    RECT 36.4000 90.3000 37.2000 90.4000 ;
	    RECT -1.9000 89.7000 37.2000 90.3000 ;
	    RECT 36.4000 89.6000 37.2000 89.7000 ;
      END
   END sr[3]
   PIN sr[4]
      PORT
         LAYER metal1 ;
	    RECT 6.0000 111.8000 6.8000 119.8000 ;
	    RECT 6.0000 109.6000 6.6000 111.8000 ;
	    RECT 6.0000 102.2000 6.8000 109.6000 ;
         LAYER metal2 ;
	    RECT 6.0000 109.6000 6.8000 110.4000 ;
	    RECT 6.1000 108.4000 6.7000 109.6000 ;
	    RECT 6.0000 107.6000 6.8000 108.4000 ;
         LAYER metal3 ;
	    RECT 6.0000 110.3000 6.8000 110.4000 ;
	    RECT -1.9000 109.7000 6.8000 110.3000 ;
	    RECT 6.0000 109.6000 6.8000 109.7000 ;
      END
   END sr[4]
   PIN sr[5]
      PORT
         LAYER metal1 ;
	    RECT 1.2000 111.8000 2.0000 119.8000 ;
	    RECT 1.2000 109.6000 1.8000 111.8000 ;
	    RECT 1.2000 102.2000 2.0000 109.6000 ;
         LAYER metal2 ;
	    RECT 1.2000 113.6000 2.0000 114.4000 ;
         LAYER metal3 ;
	    RECT 1.2000 114.3000 2.0000 114.4000 ;
	    RECT -1.9000 113.7000 2.0000 114.3000 ;
	    RECT 1.2000 113.6000 2.0000 113.7000 ;
      END
   END sr[5]
   PIN sr[6]
      PORT
         LAYER metal1 ;
	    RECT 1.2000 52.4000 2.0000 59.8000 ;
	    RECT 1.2000 50.2000 1.8000 52.4000 ;
	    RECT 1.2000 42.2000 2.0000 50.2000 ;
         LAYER metal2 ;
	    RECT 1.2000 53.6000 2.0000 54.4000 ;
         LAYER metal3 ;
	    RECT 1.2000 54.3000 2.0000 54.4000 ;
	    RECT -1.9000 53.7000 2.0000 54.3000 ;
	    RECT 1.2000 53.6000 2.0000 53.7000 ;
      END
   END sr[6]
   PIN sr[7]
      PORT
         LAYER metal1 ;
	    RECT 6.0000 52.4000 6.8000 59.8000 ;
	    RECT 6.0000 50.2000 6.6000 52.4000 ;
	    RECT 6.0000 42.2000 6.8000 50.2000 ;
         LAYER metal2 ;
	    RECT 6.0000 49.6000 6.8000 50.4000 ;
	    RECT 6.1000 48.4000 6.7000 49.6000 ;
	    RECT 6.0000 47.6000 6.8000 48.4000 ;
         LAYER metal3 ;
	    RECT 6.0000 50.3000 6.8000 50.4000 ;
	    RECT -1.9000 49.7000 6.8000 50.3000 ;
	    RECT 6.0000 49.6000 6.8000 49.7000 ;
      END
   END sr[7]
   OBS
         LAYER metal1 ;
	    RECT 4.4000 192.4000 5.2000 199.8000 ;
	    RECT 3.0000 191.8000 5.2000 192.4000 ;
	    RECT 7.6000 192.0000 8.4000 199.8000 ;
	    RECT 10.8000 195.2000 11.6000 199.8000 ;
	    RECT 3.0000 191.2000 3.6000 191.8000 ;
	    RECT 2.4000 190.4000 3.6000 191.2000 ;
	    RECT 7.4000 191.2000 8.4000 192.0000 ;
	    RECT 9.0000 194.6000 11.6000 195.2000 ;
	    RECT 9.0000 193.0000 9.6000 194.6000 ;
	    RECT 14.0000 194.4000 14.8000 199.8000 ;
	    RECT 17.2000 197.0000 18.0000 199.8000 ;
	    RECT 18.8000 197.0000 19.6000 199.8000 ;
	    RECT 20.4000 197.0000 21.2000 199.8000 ;
	    RECT 15.4000 194.4000 19.6000 195.2000 ;
	    RECT 12.2000 193.6000 14.8000 194.4000 ;
	    RECT 22.0000 193.6000 22.8000 199.8000 ;
	    RECT 25.2000 195.0000 26.0000 199.8000 ;
	    RECT 28.4000 195.0000 29.2000 199.8000 ;
	    RECT 30.0000 197.0000 30.8000 199.8000 ;
	    RECT 31.6000 197.0000 32.4000 199.8000 ;
	    RECT 34.8000 195.2000 35.6000 199.8000 ;
	    RECT 38.0000 196.4000 38.8000 199.8000 ;
	    RECT 38.0000 195.8000 39.0000 196.4000 ;
	    RECT 38.4000 195.2000 39.0000 195.8000 ;
	    RECT 33.6000 194.4000 37.8000 195.2000 ;
	    RECT 38.4000 194.6000 40.4000 195.2000 ;
	    RECT 25.2000 193.6000 27.8000 194.4000 ;
	    RECT 28.4000 193.8000 34.2000 194.4000 ;
	    RECT 37.2000 194.0000 37.8000 194.4000 ;
	    RECT 17.2000 193.0000 18.0000 193.2000 ;
	    RECT 9.0000 192.4000 18.0000 193.0000 ;
	    RECT 20.4000 193.0000 21.2000 193.2000 ;
	    RECT 28.4000 193.0000 29.0000 193.8000 ;
	    RECT 34.8000 193.2000 36.2000 193.8000 ;
	    RECT 37.2000 193.2000 38.8000 194.0000 ;
	    RECT 20.4000 192.4000 29.0000 193.0000 ;
	    RECT 30.0000 193.0000 36.2000 193.2000 ;
	    RECT 30.0000 192.6000 35.4000 193.0000 ;
	    RECT 30.0000 192.4000 30.8000 192.6000 ;
	    RECT 3.0000 187.4000 3.6000 190.4000 ;
	    RECT 4.4000 190.3000 5.2000 190.4000 ;
	    RECT 7.4000 190.3000 8.2000 191.2000 ;
	    RECT 9.0000 190.6000 9.6000 192.4000 ;
	    RECT 4.4000 189.7000 8.2000 190.3000 ;
	    RECT 4.4000 188.8000 5.2000 189.7000 ;
	    RECT 3.0000 186.8000 5.2000 187.4000 ;
	    RECT 4.4000 182.2000 5.2000 186.8000 ;
	    RECT 7.4000 186.8000 8.2000 189.7000 ;
	    RECT 8.8000 190.0000 9.6000 190.6000 ;
	    RECT 15.6000 190.0000 39.0000 190.6000 ;
	    RECT 8.8000 188.0000 9.4000 190.0000 ;
	    RECT 15.6000 189.4000 16.4000 190.0000 ;
	    RECT 33.2000 189.6000 34.0000 190.0000 ;
	    RECT 36.4000 189.6000 37.2000 190.0000 ;
	    RECT 38.2000 189.8000 39.0000 190.0000 ;
	    RECT 10.0000 188.6000 13.8000 189.4000 ;
	    RECT 8.8000 187.4000 10.0000 188.0000 ;
	    RECT 6.0000 186.3000 6.8000 186.4000 ;
	    RECT 7.4000 186.3000 8.4000 186.8000 ;
	    RECT 6.0000 185.7000 8.4000 186.3000 ;
	    RECT 6.0000 185.6000 6.8000 185.7000 ;
	    RECT 7.6000 182.2000 8.4000 185.7000 ;
	    RECT 9.2000 182.2000 10.0000 187.4000 ;
	    RECT 13.0000 187.4000 13.8000 188.6000 ;
	    RECT 13.0000 186.8000 14.8000 187.4000 ;
	    RECT 14.0000 186.2000 14.8000 186.8000 ;
	    RECT 18.8000 186.4000 19.6000 189.2000 ;
	    RECT 22.0000 188.6000 25.2000 189.4000 ;
	    RECT 29.0000 188.6000 31.0000 189.4000 ;
	    RECT 39.6000 189.0000 40.4000 194.6000 ;
	    RECT 44.4000 192.4000 45.2000 199.8000 ;
	    RECT 43.0000 191.8000 45.2000 192.4000 ;
	    RECT 52.4000 192.0000 53.2000 199.8000 ;
	    RECT 55.6000 195.2000 56.4000 199.8000 ;
	    RECT 43.0000 191.2000 43.6000 191.8000 ;
	    RECT 42.4000 190.4000 43.6000 191.2000 ;
	    RECT 52.2000 191.2000 53.2000 192.0000 ;
	    RECT 53.8000 194.6000 56.4000 195.2000 ;
	    RECT 53.8000 193.0000 54.4000 194.6000 ;
	    RECT 58.8000 194.4000 59.6000 199.8000 ;
	    RECT 62.0000 197.0000 62.8000 199.8000 ;
	    RECT 63.6000 197.0000 64.4000 199.8000 ;
	    RECT 65.2000 197.0000 66.0000 199.8000 ;
	    RECT 60.2000 194.4000 64.4000 195.2000 ;
	    RECT 57.0000 193.6000 59.6000 194.4000 ;
	    RECT 66.8000 193.6000 67.6000 199.8000 ;
	    RECT 70.0000 195.0000 70.8000 199.8000 ;
	    RECT 73.2000 195.0000 74.0000 199.8000 ;
	    RECT 74.8000 197.0000 75.6000 199.8000 ;
	    RECT 76.4000 197.0000 77.2000 199.8000 ;
	    RECT 79.6000 195.2000 80.4000 199.8000 ;
	    RECT 82.8000 196.4000 83.6000 199.8000 ;
	    RECT 82.8000 195.8000 83.8000 196.4000 ;
	    RECT 83.2000 195.2000 83.8000 195.8000 ;
	    RECT 78.4000 194.4000 82.6000 195.2000 ;
	    RECT 83.2000 194.6000 85.2000 195.2000 ;
	    RECT 70.0000 193.6000 72.6000 194.4000 ;
	    RECT 73.2000 193.8000 79.0000 194.4000 ;
	    RECT 82.0000 194.0000 82.6000 194.4000 ;
	    RECT 62.0000 193.0000 62.8000 193.2000 ;
	    RECT 53.8000 192.4000 62.8000 193.0000 ;
	    RECT 65.2000 193.0000 66.0000 193.2000 ;
	    RECT 73.2000 193.0000 73.8000 193.8000 ;
	    RECT 79.6000 193.2000 81.0000 193.8000 ;
	    RECT 82.0000 193.2000 83.6000 194.0000 ;
	    RECT 65.2000 192.4000 73.8000 193.0000 ;
	    RECT 74.8000 193.0000 81.0000 193.2000 ;
	    RECT 74.8000 192.6000 80.2000 193.0000 ;
	    RECT 74.8000 192.4000 75.6000 192.6000 ;
	    RECT 21.6000 187.8000 22.4000 188.0000 ;
	    RECT 21.6000 187.2000 26.0000 187.8000 ;
	    RECT 25.2000 187.0000 26.0000 187.2000 ;
	    RECT 26.8000 186.8000 27.6000 188.4000 ;
	    RECT 14.0000 185.4000 16.4000 186.2000 ;
	    RECT 18.8000 185.6000 19.8000 186.4000 ;
	    RECT 22.8000 185.6000 24.4000 186.4000 ;
	    RECT 25.2000 186.2000 26.0000 186.4000 ;
	    RECT 29.0000 186.2000 29.8000 188.6000 ;
	    RECT 31.6000 188.2000 40.4000 189.0000 ;
	    RECT 35.0000 186.8000 38.0000 187.6000 ;
	    RECT 35.0000 186.2000 35.8000 186.8000 ;
	    RECT 25.2000 185.6000 29.8000 186.2000 ;
	    RECT 15.6000 182.2000 16.4000 185.4000 ;
	    RECT 33.2000 185.4000 35.8000 186.2000 ;
	    RECT 17.2000 182.2000 18.0000 185.0000 ;
	    RECT 18.8000 182.2000 19.6000 185.0000 ;
	    RECT 20.4000 182.2000 21.2000 185.0000 ;
	    RECT 22.0000 182.2000 22.8000 185.0000 ;
	    RECT 25.2000 182.2000 26.0000 185.0000 ;
	    RECT 28.4000 182.2000 29.2000 185.0000 ;
	    RECT 30.0000 182.2000 30.8000 185.0000 ;
	    RECT 31.6000 182.2000 32.4000 185.0000 ;
	    RECT 33.2000 182.2000 34.0000 185.4000 ;
	    RECT 39.6000 182.2000 40.4000 188.2000 ;
	    RECT 43.0000 187.4000 43.6000 190.4000 ;
	    RECT 44.4000 190.3000 45.2000 190.4000 ;
	    RECT 52.2000 190.3000 53.0000 191.2000 ;
	    RECT 53.8000 190.6000 54.4000 192.4000 ;
	    RECT 44.4000 189.7000 53.0000 190.3000 ;
	    RECT 44.4000 188.8000 45.2000 189.7000 ;
	    RECT 43.0000 186.8000 45.2000 187.4000 ;
	    RECT 44.4000 182.2000 45.2000 186.8000 ;
	    RECT 52.2000 186.8000 53.0000 189.7000 ;
	    RECT 53.6000 190.0000 54.4000 190.6000 ;
	    RECT 60.4000 190.0000 83.8000 190.6000 ;
	    RECT 53.6000 188.0000 54.2000 190.0000 ;
	    RECT 60.4000 189.4000 61.2000 190.0000 ;
	    RECT 78.0000 189.6000 78.8000 190.0000 ;
	    RECT 81.2000 189.6000 82.0000 190.0000 ;
	    RECT 83.0000 189.8000 83.8000 190.0000 ;
	    RECT 54.8000 188.6000 58.6000 189.4000 ;
	    RECT 53.6000 187.4000 54.8000 188.0000 ;
	    RECT 52.2000 186.0000 53.2000 186.8000 ;
	    RECT 52.4000 182.2000 53.2000 186.0000 ;
	    RECT 54.0000 182.2000 54.8000 187.4000 ;
	    RECT 57.8000 187.4000 58.6000 188.6000 ;
	    RECT 57.8000 186.8000 59.6000 187.4000 ;
	    RECT 58.8000 186.2000 59.6000 186.8000 ;
	    RECT 63.6000 186.4000 64.4000 189.2000 ;
	    RECT 66.8000 188.6000 70.0000 189.4000 ;
	    RECT 73.8000 188.6000 75.8000 189.4000 ;
	    RECT 84.4000 189.0000 85.2000 194.6000 ;
	    RECT 89.2000 192.4000 90.0000 199.8000 ;
	    RECT 87.8000 191.8000 90.0000 192.4000 ;
	    RECT 90.8000 192.4000 91.6000 199.8000 ;
	    RECT 95.6000 192.4000 96.4000 199.8000 ;
	    RECT 90.8000 191.8000 93.0000 192.4000 ;
	    RECT 95.6000 191.8000 97.8000 192.4000 ;
	    RECT 87.8000 191.2000 88.4000 191.8000 ;
	    RECT 87.2000 190.4000 88.4000 191.2000 ;
	    RECT 92.4000 191.2000 93.0000 191.8000 ;
	    RECT 97.2000 191.2000 97.8000 191.8000 ;
	    RECT 92.4000 190.4000 93.6000 191.2000 ;
	    RECT 97.2000 190.4000 98.4000 191.2000 ;
	    RECT 66.4000 187.8000 67.2000 188.0000 ;
	    RECT 66.4000 187.2000 70.8000 187.8000 ;
	    RECT 70.0000 187.0000 70.8000 187.2000 ;
	    RECT 71.6000 186.8000 72.4000 188.4000 ;
	    RECT 58.8000 185.4000 61.2000 186.2000 ;
	    RECT 63.6000 185.6000 64.6000 186.4000 ;
	    RECT 67.6000 185.6000 69.2000 186.4000 ;
	    RECT 70.0000 186.2000 70.8000 186.4000 ;
	    RECT 73.8000 186.2000 74.6000 188.6000 ;
	    RECT 76.4000 188.2000 85.2000 189.0000 ;
	    RECT 79.8000 186.8000 82.8000 187.6000 ;
	    RECT 79.8000 186.2000 80.6000 186.8000 ;
	    RECT 70.0000 185.6000 74.6000 186.2000 ;
	    RECT 60.4000 182.2000 61.2000 185.4000 ;
	    RECT 78.0000 185.4000 80.6000 186.2000 ;
	    RECT 62.0000 182.2000 62.8000 185.0000 ;
	    RECT 63.6000 182.2000 64.4000 185.0000 ;
	    RECT 65.2000 182.2000 66.0000 185.0000 ;
	    RECT 66.8000 182.2000 67.6000 185.0000 ;
	    RECT 70.0000 182.2000 70.8000 185.0000 ;
	    RECT 73.2000 182.2000 74.0000 185.0000 ;
	    RECT 74.8000 182.2000 75.6000 185.0000 ;
	    RECT 76.4000 182.2000 77.2000 185.0000 ;
	    RECT 78.0000 182.2000 78.8000 185.4000 ;
	    RECT 84.4000 182.2000 85.2000 188.2000 ;
	    RECT 87.8000 187.4000 88.4000 190.4000 ;
	    RECT 89.2000 188.8000 90.0000 190.4000 ;
	    RECT 90.8000 188.8000 91.6000 190.4000 ;
	    RECT 92.4000 187.4000 93.0000 190.4000 ;
	    RECT 95.6000 188.8000 96.4000 190.4000 ;
	    RECT 97.2000 187.4000 97.8000 190.4000 ;
	    RECT 87.8000 186.8000 90.0000 187.4000 ;
	    RECT 89.2000 182.2000 90.0000 186.8000 ;
	    RECT 90.8000 186.8000 93.0000 187.4000 ;
	    RECT 95.6000 186.8000 97.8000 187.4000 ;
	    RECT 102.0000 190.3000 102.8000 199.8000 ;
	    RECT 103.6000 192.4000 104.4000 199.8000 ;
	    RECT 106.8000 192.4000 107.6000 199.8000 ;
	    RECT 103.6000 191.8000 107.6000 192.4000 ;
	    RECT 108.4000 191.8000 109.2000 199.8000 ;
	    RECT 110.6000 192.6000 111.4000 199.8000 ;
	    RECT 116.4000 196.4000 117.2000 199.8000 ;
	    RECT 116.2000 195.8000 117.2000 196.4000 ;
	    RECT 116.2000 195.2000 116.8000 195.8000 ;
	    RECT 119.6000 195.2000 120.4000 199.8000 ;
	    RECT 122.8000 197.0000 123.6000 199.8000 ;
	    RECT 124.4000 197.0000 125.2000 199.8000 ;
	    RECT 114.8000 194.6000 116.8000 195.2000 ;
	    RECT 110.6000 191.8000 112.4000 192.6000 ;
	    RECT 104.4000 190.4000 105.2000 190.8000 ;
	    RECT 108.4000 190.4000 109.0000 191.8000 ;
	    RECT 103.6000 190.3000 105.2000 190.4000 ;
	    RECT 102.0000 189.8000 105.2000 190.3000 ;
	    RECT 106.8000 189.8000 109.2000 190.4000 ;
	    RECT 102.0000 189.7000 104.4000 189.8000 ;
	    RECT 90.8000 182.2000 91.6000 186.8000 ;
	    RECT 95.6000 182.2000 96.4000 186.8000 ;
	    RECT 100.4000 184.8000 101.2000 186.4000 ;
	    RECT 102.0000 182.2000 102.8000 189.7000 ;
	    RECT 103.6000 189.6000 104.4000 189.7000 ;
	    RECT 105.2000 187.6000 106.0000 189.2000 ;
	    RECT 106.8000 188.3000 107.4000 189.8000 ;
	    RECT 108.4000 189.6000 109.2000 189.8000 ;
	    RECT 110.0000 189.6000 110.8000 191.2000 ;
	    RECT 111.6000 188.4000 112.2000 191.8000 ;
	    RECT 114.8000 189.0000 115.6000 194.6000 ;
	    RECT 117.4000 194.4000 121.6000 195.2000 ;
	    RECT 126.0000 195.0000 126.8000 199.8000 ;
	    RECT 129.2000 195.0000 130.0000 199.8000 ;
	    RECT 117.4000 194.0000 118.0000 194.4000 ;
	    RECT 116.4000 193.2000 118.0000 194.0000 ;
	    RECT 121.0000 193.8000 126.8000 194.4000 ;
	    RECT 119.0000 193.2000 120.4000 193.8000 ;
	    RECT 119.0000 193.0000 125.2000 193.2000 ;
	    RECT 119.8000 192.6000 125.2000 193.0000 ;
	    RECT 124.4000 192.4000 125.2000 192.6000 ;
	    RECT 126.2000 193.0000 126.8000 193.8000 ;
	    RECT 127.4000 193.6000 130.0000 194.4000 ;
	    RECT 132.4000 193.6000 133.2000 199.8000 ;
	    RECT 134.0000 197.0000 134.8000 199.8000 ;
	    RECT 135.6000 197.0000 136.4000 199.8000 ;
	    RECT 137.2000 197.0000 138.0000 199.8000 ;
	    RECT 135.6000 194.4000 139.8000 195.2000 ;
	    RECT 140.4000 194.4000 141.2000 199.8000 ;
	    RECT 143.6000 195.2000 144.4000 199.8000 ;
	    RECT 143.6000 194.6000 146.2000 195.2000 ;
	    RECT 140.4000 193.6000 143.0000 194.4000 ;
	    RECT 134.0000 193.0000 134.8000 193.2000 ;
	    RECT 126.2000 192.4000 134.8000 193.0000 ;
	    RECT 137.2000 193.0000 138.0000 193.2000 ;
	    RECT 145.6000 193.0000 146.2000 194.6000 ;
	    RECT 137.2000 192.4000 146.2000 193.0000 ;
	    RECT 145.6000 190.6000 146.2000 192.4000 ;
	    RECT 146.8000 192.0000 147.6000 199.8000 ;
	    RECT 151.6000 195.8000 152.4000 199.8000 ;
	    RECT 151.8000 195.6000 152.4000 195.8000 ;
	    RECT 154.8000 195.8000 155.6000 199.8000 ;
	    RECT 154.8000 195.6000 155.4000 195.8000 ;
	    RECT 151.8000 195.0000 155.4000 195.6000 ;
	    RECT 153.2000 192.8000 154.0000 194.4000 ;
	    RECT 154.8000 192.4000 155.4000 195.0000 ;
	    RECT 164.4000 192.4000 165.2000 199.8000 ;
	    RECT 146.8000 191.2000 147.8000 192.0000 ;
	    RECT 116.2000 190.0000 139.6000 190.6000 ;
	    RECT 145.6000 190.0000 146.4000 190.6000 ;
	    RECT 116.2000 189.8000 117.0000 190.0000 ;
	    RECT 118.0000 189.6000 118.8000 190.0000 ;
	    RECT 121.2000 189.6000 122.0000 190.0000 ;
	    RECT 138.8000 189.4000 139.6000 190.0000 ;
	    RECT 108.4000 188.3000 109.2000 188.4000 ;
	    RECT 106.8000 187.7000 109.2000 188.3000 ;
	    RECT 106.8000 186.2000 107.4000 187.7000 ;
	    RECT 108.4000 187.6000 109.2000 187.7000 ;
	    RECT 111.6000 187.6000 112.4000 188.4000 ;
	    RECT 114.8000 188.2000 123.6000 189.0000 ;
	    RECT 124.2000 188.6000 126.2000 189.4000 ;
	    RECT 130.0000 188.6000 133.2000 189.4000 ;
	    RECT 108.4000 186.3000 109.2000 186.4000 ;
	    RECT 111.6000 186.3000 112.2000 187.6000 ;
	    RECT 106.8000 182.2000 107.6000 186.2000 ;
	    RECT 108.4000 185.7000 112.3000 186.3000 ;
	    RECT 108.4000 185.6000 109.2000 185.7000 ;
	    RECT 108.2000 184.8000 109.0000 185.6000 ;
	    RECT 111.6000 184.2000 112.2000 185.7000 ;
	    RECT 113.2000 184.8000 114.0000 186.4000 ;
	    RECT 111.6000 182.2000 112.4000 184.2000 ;
	    RECT 114.8000 182.2000 115.6000 188.2000 ;
	    RECT 117.2000 186.8000 120.2000 187.6000 ;
	    RECT 119.4000 186.2000 120.2000 186.8000 ;
	    RECT 125.4000 186.2000 126.2000 188.6000 ;
	    RECT 127.6000 186.8000 128.4000 188.4000 ;
	    RECT 132.8000 187.8000 133.6000 188.0000 ;
	    RECT 129.2000 187.2000 133.6000 187.8000 ;
	    RECT 129.2000 187.0000 130.0000 187.2000 ;
	    RECT 135.6000 186.4000 136.4000 189.2000 ;
	    RECT 141.4000 188.6000 145.2000 189.4000 ;
	    RECT 141.4000 187.4000 142.2000 188.6000 ;
	    RECT 145.8000 188.0000 146.4000 190.0000 ;
	    RECT 129.2000 186.2000 130.0000 186.4000 ;
	    RECT 119.4000 185.4000 122.0000 186.2000 ;
	    RECT 125.4000 185.6000 130.0000 186.2000 ;
	    RECT 130.8000 185.6000 132.4000 186.4000 ;
	    RECT 135.4000 185.6000 136.4000 186.4000 ;
	    RECT 140.4000 186.8000 142.2000 187.4000 ;
	    RECT 145.2000 187.4000 146.4000 188.0000 ;
	    RECT 140.4000 186.2000 141.2000 186.8000 ;
	    RECT 121.2000 182.2000 122.0000 185.4000 ;
	    RECT 138.8000 185.4000 141.2000 186.2000 ;
	    RECT 122.8000 182.2000 123.6000 185.0000 ;
	    RECT 124.4000 182.2000 125.2000 185.0000 ;
	    RECT 126.0000 182.2000 126.8000 185.0000 ;
	    RECT 129.2000 182.2000 130.0000 185.0000 ;
	    RECT 132.4000 182.2000 133.2000 185.0000 ;
	    RECT 134.0000 182.2000 134.8000 185.0000 ;
	    RECT 135.6000 182.2000 136.4000 185.0000 ;
	    RECT 137.2000 182.2000 138.0000 185.0000 ;
	    RECT 138.8000 182.2000 139.6000 185.4000 ;
	    RECT 145.2000 182.2000 146.0000 187.4000 ;
	    RECT 147.0000 186.8000 147.8000 191.2000 ;
	    RECT 150.0000 190.8000 150.8000 192.4000 ;
	    RECT 154.8000 191.6000 155.6000 192.4000 ;
	    RECT 163.0000 191.8000 165.2000 192.4000 ;
	    RECT 167.6000 192.0000 168.4000 199.8000 ;
	    RECT 170.8000 195.2000 171.6000 199.8000 ;
	    RECT 151.6000 189.6000 153.2000 190.4000 ;
	    RECT 154.8000 188.4000 155.4000 191.6000 ;
	    RECT 163.0000 191.2000 163.6000 191.8000 ;
	    RECT 162.4000 190.4000 163.6000 191.2000 ;
	    RECT 167.4000 191.2000 168.4000 192.0000 ;
	    RECT 169.0000 194.6000 171.6000 195.2000 ;
	    RECT 169.0000 193.0000 169.6000 194.6000 ;
	    RECT 174.0000 194.4000 174.8000 199.8000 ;
	    RECT 177.2000 197.0000 178.0000 199.8000 ;
	    RECT 178.8000 197.0000 179.6000 199.8000 ;
	    RECT 180.4000 197.0000 181.2000 199.8000 ;
	    RECT 175.4000 194.4000 179.6000 195.2000 ;
	    RECT 172.2000 193.6000 174.8000 194.4000 ;
	    RECT 182.0000 193.6000 182.8000 199.8000 ;
	    RECT 185.2000 195.0000 186.0000 199.8000 ;
	    RECT 188.4000 195.0000 189.2000 199.8000 ;
	    RECT 190.0000 197.0000 190.8000 199.8000 ;
	    RECT 191.6000 197.0000 192.4000 199.8000 ;
	    RECT 194.8000 195.2000 195.6000 199.8000 ;
	    RECT 198.0000 196.4000 198.8000 199.8000 ;
	    RECT 198.0000 195.8000 199.0000 196.4000 ;
	    RECT 198.4000 195.2000 199.0000 195.8000 ;
	    RECT 193.6000 194.4000 197.8000 195.2000 ;
	    RECT 198.4000 194.6000 200.4000 195.2000 ;
	    RECT 185.2000 193.6000 187.8000 194.4000 ;
	    RECT 188.4000 193.8000 194.2000 194.4000 ;
	    RECT 197.2000 194.0000 197.8000 194.4000 ;
	    RECT 177.2000 193.0000 178.0000 193.2000 ;
	    RECT 169.0000 192.4000 178.0000 193.0000 ;
	    RECT 180.4000 193.0000 181.2000 193.2000 ;
	    RECT 188.4000 193.0000 189.0000 193.8000 ;
	    RECT 194.8000 193.2000 196.2000 193.8000 ;
	    RECT 197.2000 193.2000 198.8000 194.0000 ;
	    RECT 180.4000 192.4000 189.0000 193.0000 ;
	    RECT 190.0000 193.0000 196.2000 193.2000 ;
	    RECT 190.0000 192.6000 195.4000 193.0000 ;
	    RECT 190.0000 192.4000 190.8000 192.6000 ;
	    RECT 153.8000 188.2000 155.4000 188.4000 ;
	    RECT 146.8000 186.0000 147.8000 186.8000 ;
	    RECT 153.6000 187.8000 155.4000 188.2000 ;
	    RECT 146.8000 182.2000 147.6000 186.0000 ;
	    RECT 153.6000 184.3000 154.4000 187.8000 ;
	    RECT 163.0000 187.4000 163.6000 190.4000 ;
	    RECT 164.4000 188.8000 165.2000 190.4000 ;
	    RECT 163.0000 186.8000 165.2000 187.4000 ;
	    RECT 159.6000 184.3000 160.4000 184.4000 ;
	    RECT 153.6000 183.7000 160.4000 184.3000 ;
	    RECT 153.6000 182.2000 154.4000 183.7000 ;
	    RECT 159.6000 183.6000 160.4000 183.7000 ;
	    RECT 164.4000 182.2000 165.2000 186.8000 ;
	    RECT 167.4000 186.8000 168.2000 191.2000 ;
	    RECT 169.0000 190.6000 169.6000 192.4000 ;
	    RECT 168.8000 190.0000 169.6000 190.6000 ;
	    RECT 175.6000 190.0000 199.0000 190.6000 ;
	    RECT 168.8000 188.0000 169.4000 190.0000 ;
	    RECT 175.6000 189.4000 176.4000 190.0000 ;
	    RECT 193.2000 189.6000 194.0000 190.0000 ;
	    RECT 194.8000 189.6000 195.6000 190.0000 ;
	    RECT 198.2000 189.8000 199.0000 190.0000 ;
	    RECT 170.0000 188.6000 173.8000 189.4000 ;
	    RECT 168.8000 187.4000 170.0000 188.0000 ;
	    RECT 167.4000 186.0000 168.4000 186.8000 ;
	    RECT 167.6000 182.2000 168.4000 186.0000 ;
	    RECT 169.2000 182.2000 170.0000 187.4000 ;
	    RECT 173.0000 187.4000 173.8000 188.6000 ;
	    RECT 173.0000 186.8000 174.8000 187.4000 ;
	    RECT 174.0000 186.2000 174.8000 186.8000 ;
	    RECT 178.8000 186.4000 179.6000 189.2000 ;
	    RECT 182.0000 188.6000 185.2000 189.4000 ;
	    RECT 189.0000 188.6000 191.0000 189.4000 ;
	    RECT 199.6000 189.0000 200.4000 194.6000 ;
	    RECT 203.8000 192.6000 204.6000 199.8000 ;
	    RECT 202.8000 191.8000 204.6000 192.6000 ;
	    RECT 206.0000 191.8000 206.8000 199.8000 ;
	    RECT 207.6000 192.4000 208.4000 199.8000 ;
	    RECT 210.8000 192.4000 211.6000 199.8000 ;
	    RECT 207.6000 191.8000 211.6000 192.4000 ;
	    RECT 181.6000 187.8000 182.4000 188.0000 ;
	    RECT 181.6000 187.2000 186.0000 187.8000 ;
	    RECT 185.2000 187.0000 186.0000 187.2000 ;
	    RECT 174.0000 185.4000 176.4000 186.2000 ;
	    RECT 178.8000 185.6000 179.8000 186.4000 ;
	    RECT 182.8000 185.6000 184.4000 186.4000 ;
	    RECT 185.2000 186.2000 186.0000 186.4000 ;
	    RECT 189.0000 186.2000 189.8000 188.6000 ;
	    RECT 191.6000 188.2000 200.4000 189.0000 ;
	    RECT 203.0000 188.4000 203.6000 191.8000 ;
	    RECT 204.4000 189.6000 205.2000 191.2000 ;
	    RECT 206.2000 190.4000 206.8000 191.8000 ;
	    RECT 210.0000 190.4000 210.8000 190.8000 ;
	    RECT 206.0000 189.8000 208.4000 190.4000 ;
	    RECT 210.0000 190.3000 211.6000 190.4000 ;
	    RECT 212.4000 190.3000 213.2000 199.8000 ;
	    RECT 218.8000 192.4000 219.6000 199.8000 ;
	    RECT 217.4000 191.8000 219.6000 192.4000 ;
	    RECT 217.4000 191.2000 218.0000 191.8000 ;
	    RECT 216.8000 190.4000 218.0000 191.2000 ;
	    RECT 210.0000 189.8000 213.2000 190.3000 ;
	    RECT 206.0000 189.6000 206.8000 189.8000 ;
	    RECT 195.0000 186.8000 198.0000 187.6000 ;
	    RECT 195.0000 186.2000 195.8000 186.8000 ;
	    RECT 185.2000 185.6000 189.8000 186.2000 ;
	    RECT 175.6000 182.2000 176.4000 185.4000 ;
	    RECT 193.2000 185.4000 195.8000 186.2000 ;
	    RECT 177.2000 182.2000 178.0000 185.0000 ;
	    RECT 178.8000 182.2000 179.6000 185.0000 ;
	    RECT 180.4000 182.2000 181.2000 185.0000 ;
	    RECT 182.0000 182.2000 182.8000 185.0000 ;
	    RECT 185.2000 182.2000 186.0000 185.0000 ;
	    RECT 188.4000 182.2000 189.2000 185.0000 ;
	    RECT 190.0000 182.2000 190.8000 185.0000 ;
	    RECT 191.6000 182.2000 192.4000 185.0000 ;
	    RECT 193.2000 182.2000 194.0000 185.4000 ;
	    RECT 199.6000 182.2000 200.4000 188.2000 ;
	    RECT 202.8000 187.6000 203.6000 188.4000 ;
	    RECT 204.4000 188.3000 205.2000 188.4000 ;
	    RECT 207.8000 188.3000 208.4000 189.8000 ;
	    RECT 210.8000 189.7000 213.2000 189.8000 ;
	    RECT 210.8000 189.6000 211.6000 189.7000 ;
	    RECT 204.4000 187.7000 208.4000 188.3000 ;
	    RECT 204.4000 187.6000 205.2000 187.7000 ;
	    RECT 203.0000 186.3000 203.6000 187.6000 ;
	    RECT 206.0000 186.3000 206.8000 186.4000 ;
	    RECT 202.9000 185.7000 206.8000 186.3000 ;
	    RECT 207.8000 186.2000 208.4000 187.7000 ;
	    RECT 209.2000 187.6000 210.0000 189.2000 ;
	    RECT 203.0000 184.2000 203.6000 185.7000 ;
	    RECT 206.0000 185.6000 206.8000 185.7000 ;
	    RECT 206.2000 184.8000 207.0000 185.6000 ;
	    RECT 202.8000 182.2000 203.6000 184.2000 ;
	    RECT 207.6000 182.2000 208.4000 186.2000 ;
	    RECT 212.4000 182.2000 213.2000 189.7000 ;
	    RECT 217.4000 187.4000 218.0000 190.4000 ;
	    RECT 218.8000 188.8000 219.6000 190.4000 ;
	    RECT 217.4000 186.8000 219.6000 187.4000 ;
	    RECT 214.0000 184.8000 214.8000 186.4000 ;
	    RECT 218.8000 182.2000 219.6000 186.8000 ;
	    RECT 220.4000 182.2000 221.2000 199.8000 ;
	    RECT 4.4000 175.2000 5.2000 179.8000 ;
	    RECT 6.0000 175.6000 6.8000 177.2000 ;
	    RECT 3.0000 174.6000 5.2000 175.2000 ;
	    RECT 3.0000 171.6000 3.6000 174.6000 ;
	    RECT 4.4000 171.6000 5.2000 173.2000 ;
	    RECT 7.6000 172.3000 8.4000 179.8000 ;
	    RECT 13.0000 178.4000 13.8000 179.0000 ;
	    RECT 13.0000 177.6000 14.8000 178.4000 ;
	    RECT 13.0000 176.0000 13.8000 177.6000 ;
	    RECT 17.2000 177.0000 18.0000 179.0000 ;
	    RECT 12.2000 175.4000 13.8000 176.0000 ;
	    RECT 12.2000 175.0000 13.0000 175.4000 ;
	    RECT 12.2000 174.4000 12.8000 175.0000 ;
	    RECT 17.4000 174.8000 18.0000 177.0000 ;
	    RECT 20.4000 176.0000 21.2000 179.8000 ;
	    RECT 10.8000 173.6000 12.8000 174.4000 ;
	    RECT 13.8000 174.2000 18.0000 174.8000 ;
	    RECT 20.2000 175.2000 21.2000 176.0000 ;
	    RECT 13.8000 173.8000 14.8000 174.2000 ;
	    RECT 10.8000 172.3000 11.6000 172.4000 ;
	    RECT 7.6000 171.7000 11.6000 172.3000 ;
	    RECT 2.4000 170.8000 3.6000 171.6000 ;
	    RECT 3.0000 170.2000 3.6000 170.8000 ;
	    RECT 3.0000 169.6000 5.2000 170.2000 ;
	    RECT 4.4000 162.2000 5.2000 169.6000 ;
	    RECT 7.6000 162.2000 8.4000 171.7000 ;
	    RECT 10.8000 170.8000 11.6000 171.7000 ;
	    RECT 12.2000 169.8000 12.8000 173.6000 ;
	    RECT 13.4000 173.0000 14.8000 173.8000 ;
	    RECT 14.2000 171.0000 14.8000 173.0000 ;
	    RECT 15.6000 171.6000 16.4000 173.2000 ;
	    RECT 17.2000 171.6000 18.0000 173.2000 ;
	    RECT 14.2000 170.4000 18.0000 171.0000 ;
	    RECT 12.2000 169.2000 13.8000 169.8000 ;
	    RECT 13.0000 162.2000 13.8000 169.2000 ;
	    RECT 17.4000 167.0000 18.0000 170.4000 ;
	    RECT 20.2000 170.8000 21.0000 175.2000 ;
	    RECT 22.0000 174.6000 22.8000 179.8000 ;
	    RECT 28.4000 176.6000 29.2000 179.8000 ;
	    RECT 30.0000 177.0000 30.8000 179.8000 ;
	    RECT 31.6000 177.0000 32.4000 179.8000 ;
	    RECT 33.2000 177.0000 34.0000 179.8000 ;
	    RECT 34.8000 177.0000 35.6000 179.8000 ;
	    RECT 38.0000 177.0000 38.8000 179.8000 ;
	    RECT 41.2000 177.0000 42.0000 179.8000 ;
	    RECT 42.8000 177.0000 43.6000 179.8000 ;
	    RECT 44.4000 177.0000 45.2000 179.8000 ;
	    RECT 26.8000 175.8000 29.2000 176.6000 ;
	    RECT 46.0000 176.6000 46.8000 179.8000 ;
	    RECT 26.8000 175.2000 27.6000 175.8000 ;
	    RECT 21.6000 174.0000 22.8000 174.6000 ;
	    RECT 25.8000 174.6000 27.6000 175.2000 ;
	    RECT 31.6000 175.6000 32.6000 176.4000 ;
	    RECT 35.6000 175.6000 37.2000 176.4000 ;
	    RECT 38.0000 175.8000 42.6000 176.4000 ;
	    RECT 46.0000 175.8000 48.6000 176.6000 ;
	    RECT 38.0000 175.6000 38.8000 175.8000 ;
	    RECT 21.6000 172.0000 22.2000 174.0000 ;
	    RECT 25.8000 173.4000 26.6000 174.6000 ;
	    RECT 22.8000 172.6000 26.6000 173.4000 ;
	    RECT 31.6000 172.8000 32.4000 175.6000 ;
	    RECT 38.0000 174.8000 38.8000 175.0000 ;
	    RECT 34.4000 174.2000 38.8000 174.8000 ;
	    RECT 34.4000 174.0000 35.2000 174.2000 ;
	    RECT 39.6000 173.6000 40.4000 175.2000 ;
	    RECT 41.8000 173.4000 42.6000 175.8000 ;
	    RECT 47.8000 175.2000 48.6000 175.8000 ;
	    RECT 47.8000 174.4000 50.8000 175.2000 ;
	    RECT 52.4000 173.8000 53.2000 179.8000 ;
	    RECT 54.0000 175.6000 54.8000 177.2000 ;
	    RECT 34.8000 172.6000 38.0000 173.4000 ;
	    RECT 41.8000 172.6000 43.8000 173.4000 ;
	    RECT 44.4000 173.0000 53.2000 173.8000 ;
	    RECT 28.4000 172.0000 29.2000 172.6000 ;
	    RECT 39.6000 172.0000 40.4000 172.4000 ;
	    RECT 46.0000 172.0000 46.8000 172.4000 ;
	    RECT 49.2000 172.0000 50.0000 172.4000 ;
	    RECT 51.0000 172.0000 51.8000 172.2000 ;
	    RECT 21.6000 171.4000 22.4000 172.0000 ;
	    RECT 28.4000 171.4000 51.8000 172.0000 ;
	    RECT 20.2000 170.0000 21.2000 170.8000 ;
	    RECT 17.2000 163.0000 18.0000 167.0000 ;
	    RECT 20.4000 162.2000 21.2000 170.0000 ;
	    RECT 21.8000 169.6000 22.4000 171.4000 ;
	    RECT 21.8000 169.0000 30.8000 169.6000 ;
	    RECT 21.8000 167.4000 22.4000 169.0000 ;
	    RECT 30.0000 168.8000 30.8000 169.0000 ;
	    RECT 33.2000 169.0000 41.8000 169.6000 ;
	    RECT 33.2000 168.8000 34.0000 169.0000 ;
	    RECT 25.0000 167.6000 27.6000 168.4000 ;
	    RECT 21.8000 166.8000 24.4000 167.4000 ;
	    RECT 23.6000 162.2000 24.4000 166.8000 ;
	    RECT 26.8000 162.2000 27.6000 167.6000 ;
	    RECT 28.2000 166.8000 32.4000 167.6000 ;
	    RECT 30.0000 162.2000 30.8000 165.0000 ;
	    RECT 31.6000 162.2000 32.4000 165.0000 ;
	    RECT 33.2000 162.2000 34.0000 165.0000 ;
	    RECT 34.8000 162.2000 35.6000 168.4000 ;
	    RECT 38.0000 167.6000 40.6000 168.4000 ;
	    RECT 41.2000 168.2000 41.8000 169.0000 ;
	    RECT 42.8000 169.4000 43.6000 169.6000 ;
	    RECT 42.8000 169.0000 48.2000 169.4000 ;
	    RECT 42.8000 168.8000 49.0000 169.0000 ;
	    RECT 47.6000 168.2000 49.0000 168.8000 ;
	    RECT 41.2000 167.6000 47.0000 168.2000 ;
	    RECT 50.0000 168.0000 51.6000 168.8000 ;
	    RECT 50.0000 167.6000 50.6000 168.0000 ;
	    RECT 38.0000 162.2000 38.8000 167.0000 ;
	    RECT 41.2000 162.2000 42.0000 167.0000 ;
	    RECT 46.4000 166.8000 50.6000 167.6000 ;
	    RECT 52.4000 167.4000 53.2000 173.0000 ;
	    RECT 51.2000 166.8000 53.2000 167.4000 ;
	    RECT 55.6000 172.3000 56.4000 179.8000 ;
	    RECT 57.2000 175.6000 58.0000 177.2000 ;
	    RECT 57.2000 172.3000 58.0000 172.4000 ;
	    RECT 55.6000 171.7000 58.0000 172.3000 ;
	    RECT 42.8000 162.2000 43.6000 165.0000 ;
	    RECT 44.4000 162.2000 45.2000 165.0000 ;
	    RECT 47.6000 162.2000 48.4000 166.8000 ;
	    RECT 51.2000 166.2000 51.8000 166.8000 ;
	    RECT 50.8000 165.6000 51.8000 166.2000 ;
	    RECT 50.8000 162.2000 51.6000 165.6000 ;
	    RECT 55.6000 162.2000 56.4000 171.7000 ;
	    RECT 57.2000 171.6000 58.0000 171.7000 ;
	    RECT 58.8000 172.3000 59.6000 179.8000 ;
	    RECT 69.0000 178.4000 69.8000 179.0000 ;
	    RECT 69.0000 177.6000 70.8000 178.4000 ;
	    RECT 69.0000 176.0000 69.8000 177.6000 ;
	    RECT 73.2000 177.0000 74.0000 179.0000 ;
	    RECT 68.2000 175.4000 69.8000 176.0000 ;
	    RECT 68.2000 175.0000 69.0000 175.4000 ;
	    RECT 68.2000 174.4000 68.8000 175.0000 ;
	    RECT 73.4000 174.8000 74.0000 177.0000 ;
	    RECT 66.8000 173.6000 68.8000 174.4000 ;
	    RECT 69.8000 174.2000 74.0000 174.8000 ;
	    RECT 78.0000 175.8000 78.8000 179.8000 ;
	    RECT 79.4000 176.4000 80.2000 177.2000 ;
	    RECT 69.8000 173.8000 70.8000 174.2000 ;
	    RECT 66.8000 172.3000 67.6000 172.4000 ;
	    RECT 58.8000 171.7000 67.6000 172.3000 ;
	    RECT 58.8000 162.2000 59.6000 171.7000 ;
	    RECT 66.8000 170.8000 67.6000 171.7000 ;
	    RECT 68.2000 169.8000 68.8000 173.6000 ;
	    RECT 69.4000 173.0000 70.8000 173.8000 ;
	    RECT 70.2000 171.0000 70.8000 173.0000 ;
	    RECT 71.6000 171.6000 72.4000 173.2000 ;
	    RECT 73.2000 171.6000 74.0000 173.2000 ;
	    RECT 76.4000 172.8000 77.2000 174.4000 ;
	    RECT 74.8000 172.2000 75.6000 172.4000 ;
	    RECT 78.0000 172.2000 78.6000 175.8000 ;
	    RECT 79.6000 175.6000 80.4000 176.4000 ;
	    RECT 81.2000 176.0000 82.0000 179.8000 ;
	    RECT 84.4000 176.0000 85.2000 179.8000 ;
	    RECT 81.2000 175.8000 85.2000 176.0000 ;
	    RECT 86.0000 175.8000 86.8000 179.8000 ;
	    RECT 89.2000 176.0000 90.0000 179.8000 ;
	    RECT 81.4000 175.4000 85.0000 175.8000 ;
	    RECT 82.0000 174.4000 82.8000 174.8000 ;
	    RECT 86.0000 174.4000 86.6000 175.8000 ;
	    RECT 89.0000 175.2000 90.0000 176.0000 ;
	    RECT 81.2000 173.8000 82.8000 174.4000 ;
	    RECT 81.2000 173.6000 82.0000 173.8000 ;
	    RECT 84.2000 173.6000 86.8000 174.4000 ;
	    RECT 79.6000 172.2000 80.4000 172.4000 ;
	    RECT 74.8000 171.6000 76.4000 172.2000 ;
	    RECT 78.0000 171.6000 80.4000 172.2000 ;
	    RECT 82.8000 171.6000 83.6000 173.2000 ;
	    RECT 75.6000 171.2000 76.4000 171.6000 ;
	    RECT 70.2000 170.4000 74.0000 171.0000 ;
	    RECT 68.2000 169.2000 69.8000 169.8000 ;
	    RECT 69.0000 162.2000 69.8000 169.2000 ;
	    RECT 73.4000 167.0000 74.0000 170.4000 ;
	    RECT 79.6000 170.2000 80.2000 171.6000 ;
	    RECT 84.2000 170.2000 84.8000 173.6000 ;
	    RECT 89.0000 170.8000 89.8000 175.2000 ;
	    RECT 90.8000 174.6000 91.6000 179.8000 ;
	    RECT 97.2000 176.6000 98.0000 179.8000 ;
	    RECT 98.8000 177.0000 99.6000 179.8000 ;
	    RECT 100.4000 177.0000 101.2000 179.8000 ;
	    RECT 102.0000 177.0000 102.8000 179.8000 ;
	    RECT 103.6000 177.0000 104.4000 179.8000 ;
	    RECT 106.8000 177.0000 107.6000 179.8000 ;
	    RECT 110.0000 177.0000 110.8000 179.8000 ;
	    RECT 111.6000 177.0000 112.4000 179.8000 ;
	    RECT 113.2000 177.0000 114.0000 179.8000 ;
	    RECT 95.6000 175.8000 98.0000 176.6000 ;
	    RECT 114.8000 176.6000 115.6000 179.8000 ;
	    RECT 95.6000 175.2000 96.4000 175.8000 ;
	    RECT 90.4000 174.0000 91.6000 174.6000 ;
	    RECT 94.6000 174.6000 96.4000 175.2000 ;
	    RECT 100.4000 175.6000 101.4000 176.4000 ;
	    RECT 104.4000 175.6000 106.0000 176.4000 ;
	    RECT 106.8000 175.8000 111.4000 176.4000 ;
	    RECT 114.8000 175.8000 117.4000 176.6000 ;
	    RECT 106.8000 175.6000 107.6000 175.8000 ;
	    RECT 90.4000 172.0000 91.0000 174.0000 ;
	    RECT 94.6000 173.4000 95.4000 174.6000 ;
	    RECT 91.6000 172.6000 95.4000 173.4000 ;
	    RECT 100.4000 172.8000 101.2000 175.6000 ;
	    RECT 106.8000 174.8000 107.6000 175.0000 ;
	    RECT 103.2000 174.2000 107.6000 174.8000 ;
	    RECT 103.2000 174.0000 104.0000 174.2000 ;
	    RECT 108.4000 173.6000 109.2000 175.2000 ;
	    RECT 110.6000 173.4000 111.4000 175.8000 ;
	    RECT 116.6000 175.2000 117.4000 175.8000 ;
	    RECT 116.6000 174.4000 119.6000 175.2000 ;
	    RECT 121.2000 173.8000 122.0000 179.8000 ;
	    RECT 103.6000 172.6000 106.8000 173.4000 ;
	    RECT 110.6000 172.6000 112.6000 173.4000 ;
	    RECT 113.2000 173.0000 122.0000 173.8000 ;
	    RECT 97.2000 172.0000 98.0000 172.6000 ;
	    RECT 114.8000 172.0000 115.6000 172.4000 ;
	    RECT 118.0000 172.0000 118.8000 172.4000 ;
	    RECT 119.8000 172.0000 120.6000 172.2000 ;
	    RECT 90.4000 171.4000 91.2000 172.0000 ;
	    RECT 97.2000 171.4000 120.6000 172.0000 ;
	    RECT 86.0000 170.3000 86.8000 170.4000 ;
	    RECT 87.6000 170.3000 88.4000 170.4000 ;
	    RECT 86.0000 170.2000 88.4000 170.3000 ;
	    RECT 73.2000 163.0000 74.0000 167.0000 ;
	    RECT 74.8000 169.6000 78.8000 170.2000 ;
	    RECT 74.8000 162.2000 75.6000 169.6000 ;
	    RECT 78.0000 162.2000 78.8000 169.6000 ;
	    RECT 79.6000 162.2000 80.4000 170.2000 ;
	    RECT 83.8000 169.6000 84.8000 170.2000 ;
	    RECT 85.4000 169.7000 88.4000 170.2000 ;
	    RECT 89.0000 170.0000 90.0000 170.8000 ;
	    RECT 85.4000 169.6000 86.8000 169.7000 ;
	    RECT 87.6000 169.6000 88.4000 169.7000 ;
	    RECT 83.8000 162.2000 84.6000 169.6000 ;
	    RECT 85.4000 168.4000 86.0000 169.6000 ;
	    RECT 85.2000 167.6000 86.0000 168.4000 ;
	    RECT 89.2000 162.2000 90.0000 170.0000 ;
	    RECT 90.6000 169.6000 91.2000 171.4000 ;
	    RECT 90.6000 169.0000 99.6000 169.6000 ;
	    RECT 90.6000 167.4000 91.2000 169.0000 ;
	    RECT 98.8000 168.8000 99.6000 169.0000 ;
	    RECT 102.0000 169.0000 110.6000 169.6000 ;
	    RECT 102.0000 168.8000 102.8000 169.0000 ;
	    RECT 93.8000 167.6000 96.4000 168.4000 ;
	    RECT 90.6000 166.8000 93.2000 167.4000 ;
	    RECT 92.4000 162.2000 93.2000 166.8000 ;
	    RECT 95.6000 162.2000 96.4000 167.6000 ;
	    RECT 97.0000 166.8000 101.2000 167.6000 ;
	    RECT 98.8000 162.2000 99.6000 165.0000 ;
	    RECT 100.4000 162.2000 101.2000 165.0000 ;
	    RECT 102.0000 162.2000 102.8000 165.0000 ;
	    RECT 103.6000 162.2000 104.4000 168.4000 ;
	    RECT 106.8000 167.6000 109.4000 168.4000 ;
	    RECT 110.0000 168.2000 110.6000 169.0000 ;
	    RECT 111.6000 169.4000 112.4000 169.6000 ;
	    RECT 111.6000 169.0000 117.0000 169.4000 ;
	    RECT 111.6000 168.8000 117.8000 169.0000 ;
	    RECT 116.4000 168.2000 117.8000 168.8000 ;
	    RECT 110.0000 167.6000 115.8000 168.2000 ;
	    RECT 118.8000 168.0000 120.4000 168.8000 ;
	    RECT 118.8000 167.6000 119.4000 168.0000 ;
	    RECT 106.8000 162.2000 107.6000 167.0000 ;
	    RECT 110.0000 162.2000 110.8000 167.0000 ;
	    RECT 115.2000 166.8000 119.4000 167.6000 ;
	    RECT 121.2000 167.4000 122.0000 173.0000 ;
	    RECT 120.0000 166.8000 122.0000 167.4000 ;
	    RECT 122.8000 172.4000 123.6000 179.8000 ;
	    RECT 126.0000 175.2000 126.8000 179.8000 ;
	    RECT 124.6000 174.6000 126.8000 175.2000 ;
	    RECT 127.6000 177.0000 128.4000 179.0000 ;
	    RECT 131.8000 178.4000 132.6000 179.0000 ;
	    RECT 130.8000 177.6000 132.6000 178.4000 ;
	    RECT 127.6000 174.8000 128.2000 177.0000 ;
	    RECT 131.8000 176.0000 132.6000 177.6000 ;
	    RECT 131.8000 175.4000 133.4000 176.0000 ;
	    RECT 132.6000 175.0000 133.4000 175.4000 ;
	    RECT 122.8000 170.2000 123.4000 172.4000 ;
	    RECT 124.6000 171.6000 125.2000 174.6000 ;
	    RECT 127.6000 174.2000 131.8000 174.8000 ;
	    RECT 130.8000 173.8000 131.8000 174.2000 ;
	    RECT 132.8000 174.4000 133.4000 175.0000 ;
	    RECT 126.0000 171.6000 126.8000 173.2000 ;
	    RECT 127.6000 171.6000 128.4000 173.2000 ;
	    RECT 129.2000 171.6000 130.0000 173.2000 ;
	    RECT 130.8000 173.0000 132.2000 173.8000 ;
	    RECT 132.8000 173.6000 134.8000 174.4000 ;
	    RECT 124.0000 170.8000 125.2000 171.6000 ;
	    RECT 130.8000 171.0000 131.4000 173.0000 ;
	    RECT 124.6000 170.2000 125.2000 170.8000 ;
	    RECT 127.6000 170.4000 131.4000 171.0000 ;
	    RECT 111.6000 162.2000 112.4000 165.0000 ;
	    RECT 113.2000 162.2000 114.0000 165.0000 ;
	    RECT 116.4000 162.2000 117.2000 166.8000 ;
	    RECT 120.0000 166.2000 120.6000 166.8000 ;
	    RECT 119.6000 165.6000 120.6000 166.2000 ;
	    RECT 119.6000 162.2000 120.4000 165.6000 ;
	    RECT 122.8000 162.2000 123.6000 170.2000 ;
	    RECT 124.6000 169.6000 126.8000 170.2000 ;
	    RECT 126.0000 162.2000 126.8000 169.6000 ;
	    RECT 127.6000 167.0000 128.2000 170.4000 ;
	    RECT 132.8000 169.8000 133.4000 173.6000 ;
	    RECT 134.0000 172.3000 134.8000 172.4000 ;
	    RECT 135.6000 172.3000 136.4000 172.4000 ;
	    RECT 134.0000 171.7000 136.4000 172.3000 ;
	    RECT 134.0000 170.8000 134.8000 171.7000 ;
	    RECT 135.6000 171.6000 136.4000 171.7000 ;
	    RECT 131.8000 169.2000 133.4000 169.8000 ;
	    RECT 127.6000 163.0000 128.4000 167.0000 ;
	    RECT 131.8000 162.2000 132.6000 169.2000 ;
	    RECT 137.2000 162.2000 138.0000 179.8000 ;
	    RECT 138.8000 172.3000 139.6000 172.4000 ;
	    RECT 140.4000 172.3000 141.2000 179.8000 ;
	    RECT 145.2000 177.8000 146.0000 179.8000 ;
	    RECT 142.0000 175.6000 142.8000 177.2000 ;
	    RECT 143.6000 175.6000 144.4000 177.2000 ;
	    RECT 145.4000 174.4000 146.0000 177.8000 ;
	    RECT 145.2000 173.6000 146.0000 174.4000 ;
	    RECT 138.8000 171.7000 141.2000 172.3000 ;
	    RECT 138.8000 171.6000 139.6000 171.7000 ;
	    RECT 140.4000 162.2000 141.2000 171.7000 ;
	    RECT 145.4000 170.2000 146.0000 173.6000 ;
	    RECT 146.8000 172.3000 147.6000 172.4000 ;
	    RECT 148.4000 172.3000 149.2000 179.8000 ;
	    RECT 150.0000 176.3000 150.8000 177.2000 ;
	    RECT 151.6000 176.3000 152.4000 176.4000 ;
	    RECT 150.0000 175.7000 152.4000 176.3000 ;
	    RECT 158.0000 176.0000 158.8000 179.8000 ;
	    RECT 150.0000 175.6000 150.8000 175.7000 ;
	    RECT 151.6000 175.6000 152.4000 175.7000 ;
	    RECT 146.8000 171.7000 149.2000 172.3000 ;
	    RECT 146.8000 170.8000 147.6000 171.7000 ;
	    RECT 145.2000 169.4000 147.0000 170.2000 ;
	    RECT 146.2000 164.4000 147.0000 169.4000 ;
	    RECT 145.2000 163.6000 147.0000 164.4000 ;
	    RECT 146.2000 162.2000 147.0000 163.6000 ;
	    RECT 148.4000 162.2000 149.2000 171.7000 ;
	    RECT 157.8000 175.2000 158.8000 176.0000 ;
	    RECT 157.8000 170.8000 158.6000 175.2000 ;
	    RECT 159.6000 174.6000 160.4000 179.8000 ;
	    RECT 166.0000 176.6000 166.8000 179.8000 ;
	    RECT 167.6000 177.0000 168.4000 179.8000 ;
	    RECT 169.2000 177.0000 170.0000 179.8000 ;
	    RECT 170.8000 177.0000 171.6000 179.8000 ;
	    RECT 172.4000 177.0000 173.2000 179.8000 ;
	    RECT 175.6000 177.0000 176.4000 179.8000 ;
	    RECT 178.8000 177.0000 179.6000 179.8000 ;
	    RECT 180.4000 177.0000 181.2000 179.8000 ;
	    RECT 182.0000 177.0000 182.8000 179.8000 ;
	    RECT 164.4000 175.8000 166.8000 176.6000 ;
	    RECT 183.6000 176.6000 184.4000 179.8000 ;
	    RECT 164.4000 175.2000 165.2000 175.8000 ;
	    RECT 159.2000 174.0000 160.4000 174.6000 ;
	    RECT 163.4000 174.6000 165.2000 175.2000 ;
	    RECT 169.2000 175.6000 170.2000 176.4000 ;
	    RECT 173.2000 175.6000 174.8000 176.4000 ;
	    RECT 175.6000 175.8000 180.2000 176.4000 ;
	    RECT 183.6000 175.8000 186.2000 176.6000 ;
	    RECT 175.6000 175.6000 176.4000 175.8000 ;
	    RECT 159.2000 172.0000 159.8000 174.0000 ;
	    RECT 163.4000 173.4000 164.2000 174.6000 ;
	    RECT 160.4000 172.6000 164.2000 173.4000 ;
	    RECT 169.2000 172.8000 170.0000 175.6000 ;
	    RECT 175.6000 174.8000 176.4000 175.0000 ;
	    RECT 172.0000 174.2000 176.4000 174.8000 ;
	    RECT 172.0000 174.0000 172.8000 174.2000 ;
	    RECT 177.2000 173.6000 178.0000 175.2000 ;
	    RECT 179.4000 173.4000 180.2000 175.8000 ;
	    RECT 185.4000 175.2000 186.2000 175.8000 ;
	    RECT 185.4000 174.4000 188.4000 175.2000 ;
	    RECT 190.0000 173.8000 190.8000 179.8000 ;
	    RECT 172.4000 172.6000 175.6000 173.4000 ;
	    RECT 179.4000 172.6000 181.4000 173.4000 ;
	    RECT 182.0000 173.0000 190.8000 173.8000 ;
	    RECT 166.0000 172.0000 166.8000 172.6000 ;
	    RECT 183.6000 172.0000 184.4000 172.4000 ;
	    RECT 188.4000 172.2000 189.2000 172.4000 ;
	    RECT 188.4000 172.0000 189.4000 172.2000 ;
	    RECT 159.2000 171.4000 160.0000 172.0000 ;
	    RECT 166.0000 171.4000 189.4000 172.0000 ;
	    RECT 157.8000 170.0000 158.8000 170.8000 ;
	    RECT 158.0000 162.2000 158.8000 170.0000 ;
	    RECT 159.4000 169.6000 160.0000 171.4000 ;
	    RECT 159.4000 169.0000 168.4000 169.6000 ;
	    RECT 159.4000 167.4000 160.0000 169.0000 ;
	    RECT 167.6000 168.8000 168.4000 169.0000 ;
	    RECT 170.8000 169.0000 179.4000 169.6000 ;
	    RECT 170.8000 168.8000 171.6000 169.0000 ;
	    RECT 162.6000 167.6000 165.2000 168.4000 ;
	    RECT 159.4000 166.8000 162.0000 167.4000 ;
	    RECT 161.2000 162.2000 162.0000 166.8000 ;
	    RECT 164.4000 162.2000 165.2000 167.6000 ;
	    RECT 165.8000 166.8000 170.0000 167.6000 ;
	    RECT 167.6000 162.2000 168.4000 165.0000 ;
	    RECT 169.2000 162.2000 170.0000 165.0000 ;
	    RECT 170.8000 162.2000 171.6000 165.0000 ;
	    RECT 172.4000 162.2000 173.2000 168.4000 ;
	    RECT 175.6000 167.6000 178.2000 168.4000 ;
	    RECT 178.8000 168.2000 179.4000 169.0000 ;
	    RECT 180.4000 169.4000 181.2000 169.6000 ;
	    RECT 180.4000 169.0000 185.8000 169.4000 ;
	    RECT 180.4000 168.8000 186.6000 169.0000 ;
	    RECT 185.2000 168.2000 186.6000 168.8000 ;
	    RECT 178.8000 167.6000 184.6000 168.2000 ;
	    RECT 187.6000 168.0000 189.2000 168.8000 ;
	    RECT 187.6000 167.6000 188.2000 168.0000 ;
	    RECT 175.6000 162.2000 176.4000 167.0000 ;
	    RECT 178.8000 162.2000 179.6000 167.0000 ;
	    RECT 184.0000 166.8000 188.2000 167.6000 ;
	    RECT 190.0000 167.4000 190.8000 173.0000 ;
	    RECT 188.8000 166.8000 190.8000 167.4000 ;
	    RECT 191.6000 173.8000 192.4000 179.8000 ;
	    RECT 198.0000 176.6000 198.8000 179.8000 ;
	    RECT 199.6000 177.0000 200.4000 179.8000 ;
	    RECT 201.2000 177.0000 202.0000 179.8000 ;
	    RECT 202.8000 177.0000 203.6000 179.8000 ;
	    RECT 206.0000 177.0000 206.8000 179.8000 ;
	    RECT 209.2000 177.0000 210.0000 179.8000 ;
	    RECT 210.8000 177.0000 211.6000 179.8000 ;
	    RECT 212.4000 177.0000 213.2000 179.8000 ;
	    RECT 214.0000 177.0000 214.8000 179.8000 ;
	    RECT 196.2000 175.8000 198.8000 176.6000 ;
	    RECT 215.6000 176.6000 216.4000 179.8000 ;
	    RECT 202.2000 175.8000 206.8000 176.4000 ;
	    RECT 196.2000 175.2000 197.0000 175.8000 ;
	    RECT 194.0000 174.4000 197.0000 175.2000 ;
	    RECT 191.6000 173.0000 200.4000 173.8000 ;
	    RECT 202.2000 173.4000 203.0000 175.8000 ;
	    RECT 206.0000 175.6000 206.8000 175.8000 ;
	    RECT 207.6000 175.6000 209.2000 176.4000 ;
	    RECT 212.2000 175.6000 213.2000 176.4000 ;
	    RECT 215.6000 175.8000 218.0000 176.6000 ;
	    RECT 204.4000 173.6000 205.2000 175.2000 ;
	    RECT 206.0000 174.8000 206.8000 175.0000 ;
	    RECT 206.0000 174.2000 210.4000 174.8000 ;
	    RECT 209.6000 174.0000 210.4000 174.2000 ;
	    RECT 191.6000 167.4000 192.4000 173.0000 ;
	    RECT 201.0000 172.6000 203.0000 173.4000 ;
	    RECT 206.8000 172.6000 210.0000 173.4000 ;
	    RECT 212.4000 172.8000 213.2000 175.6000 ;
	    RECT 217.2000 175.2000 218.0000 175.8000 ;
	    RECT 217.2000 174.6000 219.0000 175.2000 ;
	    RECT 218.2000 173.4000 219.0000 174.6000 ;
	    RECT 222.0000 174.6000 222.8000 179.8000 ;
	    RECT 223.6000 176.0000 224.4000 179.8000 ;
	    RECT 223.6000 175.2000 224.6000 176.0000 ;
	    RECT 222.0000 174.0000 223.2000 174.6000 ;
	    RECT 218.2000 172.6000 222.0000 173.4000 ;
	    RECT 193.0000 172.0000 193.8000 172.2000 ;
	    RECT 194.8000 172.0000 195.6000 172.4000 ;
	    RECT 198.0000 172.0000 198.8000 172.4000 ;
	    RECT 215.6000 172.0000 216.4000 172.6000 ;
	    RECT 222.6000 172.0000 223.2000 174.0000 ;
	    RECT 193.0000 171.4000 216.4000 172.0000 ;
	    RECT 222.4000 171.4000 223.2000 172.0000 ;
	    RECT 222.4000 169.6000 223.0000 171.4000 ;
	    RECT 223.8000 170.8000 224.6000 175.2000 ;
	    RECT 201.2000 169.4000 202.0000 169.6000 ;
	    RECT 196.6000 169.0000 202.0000 169.4000 ;
	    RECT 195.8000 168.8000 202.0000 169.0000 ;
	    RECT 203.0000 169.0000 211.6000 169.6000 ;
	    RECT 193.2000 168.0000 194.8000 168.8000 ;
	    RECT 195.8000 168.2000 197.2000 168.8000 ;
	    RECT 203.0000 168.2000 203.6000 169.0000 ;
	    RECT 210.8000 168.8000 211.6000 169.0000 ;
	    RECT 214.0000 169.0000 223.0000 169.6000 ;
	    RECT 214.0000 168.8000 214.8000 169.0000 ;
	    RECT 194.2000 167.6000 194.8000 168.0000 ;
	    RECT 197.8000 167.6000 203.6000 168.2000 ;
	    RECT 204.2000 167.6000 206.8000 168.4000 ;
	    RECT 191.6000 166.8000 193.6000 167.4000 ;
	    RECT 194.2000 166.8000 198.4000 167.6000 ;
	    RECT 180.4000 162.2000 181.2000 165.0000 ;
	    RECT 182.0000 162.2000 182.8000 165.0000 ;
	    RECT 185.2000 162.2000 186.0000 166.8000 ;
	    RECT 188.8000 166.2000 189.4000 166.8000 ;
	    RECT 188.4000 165.6000 189.4000 166.2000 ;
	    RECT 193.0000 166.2000 193.6000 166.8000 ;
	    RECT 193.0000 165.6000 194.0000 166.2000 ;
	    RECT 188.4000 162.2000 189.2000 165.6000 ;
	    RECT 193.2000 162.2000 194.0000 165.6000 ;
	    RECT 196.4000 162.2000 197.2000 166.8000 ;
	    RECT 199.6000 162.2000 200.4000 165.0000 ;
	    RECT 201.2000 162.2000 202.0000 165.0000 ;
	    RECT 202.8000 162.2000 203.6000 167.0000 ;
	    RECT 206.0000 162.2000 206.8000 167.0000 ;
	    RECT 209.2000 162.2000 210.0000 168.4000 ;
	    RECT 217.2000 167.6000 219.8000 168.4000 ;
	    RECT 212.4000 166.8000 216.6000 167.6000 ;
	    RECT 210.8000 162.2000 211.6000 165.0000 ;
	    RECT 212.4000 162.2000 213.2000 165.0000 ;
	    RECT 214.0000 162.2000 214.8000 165.0000 ;
	    RECT 217.2000 162.2000 218.0000 167.6000 ;
	    RECT 222.4000 167.4000 223.0000 169.0000 ;
	    RECT 220.4000 166.8000 223.0000 167.4000 ;
	    RECT 223.6000 170.0000 224.6000 170.8000 ;
	    RECT 220.4000 162.2000 221.2000 166.8000 ;
	    RECT 223.6000 162.2000 224.4000 170.0000 ;
	    RECT 4.4000 152.4000 5.2000 159.8000 ;
	    RECT 3.0000 151.8000 5.2000 152.4000 ;
	    RECT 7.6000 152.0000 8.4000 159.8000 ;
	    RECT 10.8000 155.2000 11.6000 159.8000 ;
	    RECT 3.0000 151.2000 3.6000 151.8000 ;
	    RECT 2.4000 150.4000 3.6000 151.2000 ;
	    RECT 7.4000 151.2000 8.4000 152.0000 ;
	    RECT 9.0000 154.6000 11.6000 155.2000 ;
	    RECT 9.0000 153.0000 9.6000 154.6000 ;
	    RECT 14.0000 154.4000 14.8000 159.8000 ;
	    RECT 17.2000 157.0000 18.0000 159.8000 ;
	    RECT 18.8000 157.0000 19.6000 159.8000 ;
	    RECT 20.4000 157.0000 21.2000 159.8000 ;
	    RECT 15.4000 154.4000 19.6000 155.2000 ;
	    RECT 12.2000 153.6000 14.8000 154.4000 ;
	    RECT 22.0000 153.6000 22.8000 159.8000 ;
	    RECT 25.2000 155.0000 26.0000 159.8000 ;
	    RECT 28.4000 155.0000 29.2000 159.8000 ;
	    RECT 30.0000 157.0000 30.8000 159.8000 ;
	    RECT 31.6000 157.0000 32.4000 159.8000 ;
	    RECT 34.8000 155.2000 35.6000 159.8000 ;
	    RECT 38.0000 156.4000 38.8000 159.8000 ;
	    RECT 38.0000 155.8000 39.0000 156.4000 ;
	    RECT 38.4000 155.2000 39.0000 155.8000 ;
	    RECT 33.6000 154.4000 37.8000 155.2000 ;
	    RECT 38.4000 154.6000 40.4000 155.2000 ;
	    RECT 25.2000 153.6000 27.8000 154.4000 ;
	    RECT 28.4000 153.8000 34.2000 154.4000 ;
	    RECT 37.2000 154.0000 37.8000 154.4000 ;
	    RECT 17.2000 153.0000 18.0000 153.2000 ;
	    RECT 9.0000 152.4000 18.0000 153.0000 ;
	    RECT 20.4000 153.0000 21.2000 153.2000 ;
	    RECT 28.4000 153.0000 29.0000 153.8000 ;
	    RECT 34.8000 153.2000 36.2000 153.8000 ;
	    RECT 37.2000 153.2000 38.8000 154.0000 ;
	    RECT 20.4000 152.4000 29.0000 153.0000 ;
	    RECT 30.0000 153.0000 36.2000 153.2000 ;
	    RECT 30.0000 152.6000 35.4000 153.0000 ;
	    RECT 30.0000 152.4000 30.8000 152.6000 ;
	    RECT 3.0000 147.4000 3.6000 150.4000 ;
	    RECT 4.4000 150.3000 5.2000 150.4000 ;
	    RECT 7.4000 150.3000 8.2000 151.2000 ;
	    RECT 9.0000 150.6000 9.6000 152.4000 ;
	    RECT 4.4000 149.7000 8.2000 150.3000 ;
	    RECT 4.4000 148.8000 5.2000 149.7000 ;
	    RECT 3.0000 146.8000 5.2000 147.4000 ;
	    RECT 4.4000 142.2000 5.2000 146.8000 ;
	    RECT 7.4000 146.8000 8.2000 149.7000 ;
	    RECT 8.8000 150.0000 9.6000 150.6000 ;
	    RECT 15.6000 150.0000 39.0000 150.6000 ;
	    RECT 8.8000 148.0000 9.4000 150.0000 ;
	    RECT 15.6000 149.4000 16.4000 150.0000 ;
	    RECT 33.2000 149.6000 34.0000 150.0000 ;
	    RECT 36.4000 149.6000 37.2000 150.0000 ;
	    RECT 38.2000 149.8000 39.0000 150.0000 ;
	    RECT 10.0000 148.6000 13.8000 149.4000 ;
	    RECT 8.8000 147.4000 10.0000 148.0000 ;
	    RECT 6.0000 146.3000 6.8000 146.4000 ;
	    RECT 7.4000 146.3000 8.4000 146.8000 ;
	    RECT 6.0000 145.7000 8.4000 146.3000 ;
	    RECT 6.0000 145.6000 6.8000 145.7000 ;
	    RECT 7.6000 142.2000 8.4000 145.7000 ;
	    RECT 9.2000 142.2000 10.0000 147.4000 ;
	    RECT 13.0000 147.4000 13.8000 148.6000 ;
	    RECT 13.0000 146.8000 14.8000 147.4000 ;
	    RECT 14.0000 146.2000 14.8000 146.8000 ;
	    RECT 18.8000 146.4000 19.6000 149.2000 ;
	    RECT 22.0000 148.6000 25.2000 149.4000 ;
	    RECT 29.0000 148.6000 31.0000 149.4000 ;
	    RECT 39.6000 149.0000 40.4000 154.6000 ;
	    RECT 42.0000 153.6000 42.8000 154.4000 ;
	    RECT 42.0000 152.4000 42.6000 153.6000 ;
	    RECT 43.4000 152.4000 44.2000 159.8000 ;
	    RECT 41.2000 151.8000 42.6000 152.4000 ;
	    RECT 43.2000 151.8000 44.2000 152.4000 ;
	    RECT 47.6000 151.8000 48.4000 159.8000 ;
	    RECT 49.2000 152.4000 50.0000 159.8000 ;
	    RECT 52.4000 152.4000 53.2000 159.8000 ;
	    RECT 49.2000 151.8000 53.2000 152.4000 ;
	    RECT 55.6000 158.3000 56.4000 159.8000 ;
	    RECT 60.4000 158.3000 61.2000 158.4000 ;
	    RECT 55.6000 157.7000 61.2000 158.3000 ;
	    RECT 41.2000 151.6000 42.0000 151.8000 ;
	    RECT 21.6000 147.8000 22.4000 148.0000 ;
	    RECT 21.6000 147.2000 26.0000 147.8000 ;
	    RECT 25.2000 147.0000 26.0000 147.2000 ;
	    RECT 26.8000 146.8000 27.6000 148.4000 ;
	    RECT 14.0000 145.4000 16.4000 146.2000 ;
	    RECT 18.8000 145.6000 19.8000 146.4000 ;
	    RECT 22.8000 145.6000 24.4000 146.4000 ;
	    RECT 25.2000 146.2000 26.0000 146.4000 ;
	    RECT 29.0000 146.2000 29.8000 148.6000 ;
	    RECT 31.6000 148.2000 40.4000 149.0000 ;
	    RECT 43.2000 148.4000 43.8000 151.8000 ;
	    RECT 47.8000 150.4000 48.4000 151.8000 ;
	    RECT 51.6000 150.4000 52.4000 150.8000 ;
	    RECT 44.4000 148.8000 45.2000 150.4000 ;
	    RECT 47.6000 149.8000 50.0000 150.4000 ;
	    RECT 51.6000 149.8000 53.2000 150.4000 ;
	    RECT 47.6000 149.6000 48.4000 149.8000 ;
	    RECT 35.0000 146.8000 38.0000 147.6000 ;
	    RECT 35.0000 146.2000 35.8000 146.8000 ;
	    RECT 25.2000 145.6000 29.8000 146.2000 ;
	    RECT 15.6000 142.2000 16.4000 145.4000 ;
	    RECT 33.2000 145.4000 35.8000 146.2000 ;
	    RECT 17.2000 142.2000 18.0000 145.0000 ;
	    RECT 18.8000 142.2000 19.6000 145.0000 ;
	    RECT 20.4000 142.2000 21.2000 145.0000 ;
	    RECT 22.0000 142.2000 22.8000 145.0000 ;
	    RECT 25.2000 142.2000 26.0000 145.0000 ;
	    RECT 28.4000 142.2000 29.2000 145.0000 ;
	    RECT 30.0000 142.2000 30.8000 145.0000 ;
	    RECT 31.6000 142.2000 32.4000 145.0000 ;
	    RECT 33.2000 142.2000 34.0000 145.4000 ;
	    RECT 39.6000 142.2000 40.4000 148.2000 ;
	    RECT 41.2000 147.6000 43.8000 148.4000 ;
	    RECT 46.0000 148.2000 46.8000 148.4000 ;
	    RECT 45.2000 147.6000 46.8000 148.2000 ;
	    RECT 41.4000 146.2000 42.0000 147.6000 ;
	    RECT 45.2000 147.2000 46.0000 147.6000 ;
	    RECT 43.0000 146.2000 46.6000 146.6000 ;
	    RECT 41.2000 142.2000 42.0000 146.2000 ;
	    RECT 42.8000 146.0000 46.8000 146.2000 ;
	    RECT 42.8000 142.2000 43.6000 146.0000 ;
	    RECT 46.0000 142.2000 46.8000 146.0000 ;
	    RECT 47.6000 145.6000 48.4000 146.4000 ;
	    RECT 49.4000 146.2000 50.0000 149.8000 ;
	    RECT 52.4000 149.6000 53.2000 149.8000 ;
	    RECT 50.8000 148.3000 51.6000 149.2000 ;
	    RECT 55.6000 148.3000 56.4000 157.7000 ;
	    RECT 60.4000 157.6000 61.2000 157.7000 ;
	    RECT 63.6000 156.4000 64.4000 159.8000 ;
	    RECT 63.4000 155.8000 64.4000 156.4000 ;
	    RECT 63.4000 155.2000 64.0000 155.8000 ;
	    RECT 66.8000 155.2000 67.6000 159.8000 ;
	    RECT 70.0000 157.0000 70.8000 159.8000 ;
	    RECT 71.6000 157.0000 72.4000 159.8000 ;
	    RECT 50.8000 147.7000 56.4000 148.3000 ;
	    RECT 50.8000 147.6000 51.6000 147.7000 ;
	    RECT 47.8000 144.8000 48.6000 145.6000 ;
	    RECT 49.2000 142.2000 50.0000 146.2000 ;
	    RECT 54.0000 144.8000 54.8000 146.4000 ;
	    RECT 55.6000 142.2000 56.4000 147.7000 ;
	    RECT 62.0000 154.6000 64.0000 155.2000 ;
	    RECT 62.0000 149.0000 62.8000 154.6000 ;
	    RECT 64.6000 154.4000 68.8000 155.2000 ;
	    RECT 73.2000 155.0000 74.0000 159.8000 ;
	    RECT 76.4000 155.0000 77.2000 159.8000 ;
	    RECT 64.6000 154.0000 65.2000 154.4000 ;
	    RECT 63.6000 153.2000 65.2000 154.0000 ;
	    RECT 68.2000 153.8000 74.0000 154.4000 ;
	    RECT 66.2000 153.2000 67.6000 153.8000 ;
	    RECT 66.2000 153.0000 72.4000 153.2000 ;
	    RECT 67.0000 152.6000 72.4000 153.0000 ;
	    RECT 71.6000 152.4000 72.4000 152.6000 ;
	    RECT 73.4000 153.0000 74.0000 153.8000 ;
	    RECT 74.6000 153.6000 77.2000 154.4000 ;
	    RECT 79.6000 153.6000 80.4000 159.8000 ;
	    RECT 81.2000 157.0000 82.0000 159.8000 ;
	    RECT 82.8000 157.0000 83.6000 159.8000 ;
	    RECT 84.4000 157.0000 85.2000 159.8000 ;
	    RECT 82.8000 154.4000 87.0000 155.2000 ;
	    RECT 87.6000 154.4000 88.4000 159.8000 ;
	    RECT 90.8000 155.2000 91.6000 159.8000 ;
	    RECT 90.8000 154.6000 93.4000 155.2000 ;
	    RECT 87.6000 153.6000 90.2000 154.4000 ;
	    RECT 81.2000 153.0000 82.0000 153.2000 ;
	    RECT 73.4000 152.4000 82.0000 153.0000 ;
	    RECT 84.4000 153.0000 85.2000 153.2000 ;
	    RECT 92.8000 153.0000 93.4000 154.6000 ;
	    RECT 84.4000 152.4000 93.4000 153.0000 ;
	    RECT 92.8000 150.6000 93.4000 152.4000 ;
	    RECT 94.0000 154.3000 94.8000 159.8000 ;
	    RECT 98.8000 156.4000 99.6000 159.8000 ;
	    RECT 98.6000 155.8000 99.6000 156.4000 ;
	    RECT 98.6000 155.2000 99.2000 155.8000 ;
	    RECT 102.0000 155.2000 102.8000 159.8000 ;
	    RECT 105.2000 157.0000 106.0000 159.8000 ;
	    RECT 106.8000 157.0000 107.6000 159.8000 ;
	    RECT 97.2000 154.6000 99.2000 155.2000 ;
	    RECT 95.6000 154.3000 96.4000 154.4000 ;
	    RECT 94.0000 153.7000 96.4000 154.3000 ;
	    RECT 94.0000 152.0000 94.8000 153.7000 ;
	    RECT 95.6000 153.6000 96.4000 153.7000 ;
	    RECT 94.0000 151.2000 95.0000 152.0000 ;
	    RECT 63.4000 150.0000 86.8000 150.6000 ;
	    RECT 92.8000 150.0000 93.6000 150.6000 ;
	    RECT 63.4000 149.8000 64.2000 150.0000 ;
	    RECT 68.4000 149.6000 69.2000 150.0000 ;
	    RECT 86.0000 149.4000 86.8000 150.0000 ;
	    RECT 62.0000 148.2000 70.8000 149.0000 ;
	    RECT 71.4000 148.6000 73.4000 149.4000 ;
	    RECT 77.2000 148.6000 80.4000 149.4000 ;
	    RECT 62.0000 142.2000 62.8000 148.2000 ;
	    RECT 64.4000 146.8000 67.4000 147.6000 ;
	    RECT 66.6000 146.2000 67.4000 146.8000 ;
	    RECT 72.6000 146.2000 73.4000 148.6000 ;
	    RECT 74.8000 146.8000 75.6000 148.4000 ;
	    RECT 80.0000 147.8000 80.8000 148.0000 ;
	    RECT 76.4000 147.2000 80.8000 147.8000 ;
	    RECT 76.4000 147.0000 77.2000 147.2000 ;
	    RECT 82.8000 146.4000 83.6000 149.2000 ;
	    RECT 88.6000 148.6000 92.4000 149.4000 ;
	    RECT 88.6000 147.4000 89.4000 148.6000 ;
	    RECT 93.0000 148.0000 93.6000 150.0000 ;
	    RECT 76.4000 146.2000 77.2000 146.4000 ;
	    RECT 66.6000 145.4000 69.2000 146.2000 ;
	    RECT 72.6000 145.6000 77.2000 146.2000 ;
	    RECT 78.0000 145.6000 79.6000 146.4000 ;
	    RECT 82.6000 145.6000 83.6000 146.4000 ;
	    RECT 87.6000 146.8000 89.4000 147.4000 ;
	    RECT 92.4000 147.4000 93.6000 148.0000 ;
	    RECT 87.6000 146.2000 88.4000 146.8000 ;
	    RECT 68.4000 142.2000 69.2000 145.4000 ;
	    RECT 86.0000 145.4000 88.4000 146.2000 ;
	    RECT 70.0000 142.2000 70.8000 145.0000 ;
	    RECT 71.6000 142.2000 72.4000 145.0000 ;
	    RECT 73.2000 142.2000 74.0000 145.0000 ;
	    RECT 76.4000 142.2000 77.2000 145.0000 ;
	    RECT 79.6000 142.2000 80.4000 145.0000 ;
	    RECT 81.2000 142.2000 82.0000 145.0000 ;
	    RECT 82.8000 142.2000 83.6000 145.0000 ;
	    RECT 84.4000 142.2000 85.2000 145.0000 ;
	    RECT 86.0000 142.2000 86.8000 145.4000 ;
	    RECT 92.4000 142.2000 93.2000 147.4000 ;
	    RECT 94.2000 146.8000 95.0000 151.2000 ;
	    RECT 94.0000 146.0000 95.0000 146.8000 ;
	    RECT 97.2000 149.0000 98.0000 154.6000 ;
	    RECT 99.8000 154.4000 104.0000 155.2000 ;
	    RECT 108.4000 155.0000 109.2000 159.8000 ;
	    RECT 111.6000 155.0000 112.4000 159.8000 ;
	    RECT 99.8000 154.0000 100.4000 154.4000 ;
	    RECT 98.8000 153.2000 100.4000 154.0000 ;
	    RECT 103.4000 153.8000 109.2000 154.4000 ;
	    RECT 101.4000 153.2000 102.8000 153.8000 ;
	    RECT 101.4000 153.0000 107.6000 153.2000 ;
	    RECT 102.2000 152.6000 107.6000 153.0000 ;
	    RECT 106.8000 152.4000 107.6000 152.6000 ;
	    RECT 108.6000 153.0000 109.2000 153.8000 ;
	    RECT 109.8000 153.6000 112.4000 154.4000 ;
	    RECT 114.8000 153.6000 115.6000 159.8000 ;
	    RECT 116.4000 157.0000 117.2000 159.8000 ;
	    RECT 118.0000 157.0000 118.8000 159.8000 ;
	    RECT 119.6000 157.0000 120.4000 159.8000 ;
	    RECT 118.0000 154.4000 122.2000 155.2000 ;
	    RECT 122.8000 154.4000 123.6000 159.8000 ;
	    RECT 126.0000 155.2000 126.8000 159.8000 ;
	    RECT 126.0000 154.6000 128.6000 155.2000 ;
	    RECT 122.8000 153.6000 125.4000 154.4000 ;
	    RECT 116.4000 153.0000 117.2000 153.2000 ;
	    RECT 108.6000 152.4000 117.2000 153.0000 ;
	    RECT 119.6000 153.0000 120.4000 153.2000 ;
	    RECT 128.0000 153.0000 128.6000 154.6000 ;
	    RECT 119.6000 152.4000 128.6000 153.0000 ;
	    RECT 128.0000 150.6000 128.6000 152.4000 ;
	    RECT 129.2000 152.0000 130.0000 159.8000 ;
	    RECT 133.2000 153.6000 134.0000 154.4000 ;
	    RECT 133.2000 152.4000 133.8000 153.6000 ;
	    RECT 134.6000 152.4000 135.4000 159.8000 ;
	    RECT 129.2000 151.2000 130.2000 152.0000 ;
	    RECT 132.4000 151.8000 133.8000 152.4000 ;
	    RECT 134.4000 151.8000 135.4000 152.4000 ;
	    RECT 132.4000 151.6000 133.2000 151.8000 ;
	    RECT 98.6000 150.0000 122.0000 150.6000 ;
	    RECT 128.0000 150.0000 128.8000 150.6000 ;
	    RECT 98.6000 149.8000 99.4000 150.0000 ;
	    RECT 100.4000 149.6000 101.2000 150.0000 ;
	    RECT 103.6000 149.6000 104.4000 150.0000 ;
	    RECT 121.2000 149.4000 122.0000 150.0000 ;
	    RECT 97.2000 148.2000 106.0000 149.0000 ;
	    RECT 106.6000 148.6000 108.6000 149.4000 ;
	    RECT 112.4000 148.6000 115.6000 149.4000 ;
	    RECT 94.0000 142.2000 94.8000 146.0000 ;
	    RECT 97.2000 142.2000 98.0000 148.2000 ;
	    RECT 99.6000 146.8000 102.6000 147.6000 ;
	    RECT 101.8000 146.2000 102.6000 146.8000 ;
	    RECT 107.8000 146.2000 108.6000 148.6000 ;
	    RECT 110.0000 146.8000 110.8000 148.4000 ;
	    RECT 115.2000 147.8000 116.0000 148.0000 ;
	    RECT 111.6000 147.2000 116.0000 147.8000 ;
	    RECT 111.6000 147.0000 112.4000 147.2000 ;
	    RECT 118.0000 146.4000 118.8000 149.2000 ;
	    RECT 123.8000 148.6000 127.6000 149.4000 ;
	    RECT 123.8000 147.4000 124.6000 148.6000 ;
	    RECT 128.2000 148.0000 128.8000 150.0000 ;
	    RECT 111.6000 146.2000 112.4000 146.4000 ;
	    RECT 101.8000 145.4000 104.4000 146.2000 ;
	    RECT 107.8000 145.6000 112.4000 146.2000 ;
	    RECT 113.2000 145.6000 114.8000 146.4000 ;
	    RECT 117.8000 145.6000 118.8000 146.4000 ;
	    RECT 122.8000 146.8000 124.6000 147.4000 ;
	    RECT 127.6000 147.4000 128.8000 148.0000 ;
	    RECT 122.8000 146.2000 123.6000 146.8000 ;
	    RECT 103.6000 142.2000 104.4000 145.4000 ;
	    RECT 121.2000 145.4000 123.6000 146.2000 ;
	    RECT 105.2000 142.2000 106.0000 145.0000 ;
	    RECT 106.8000 142.2000 107.6000 145.0000 ;
	    RECT 108.4000 142.2000 109.2000 145.0000 ;
	    RECT 111.6000 142.2000 112.4000 145.0000 ;
	    RECT 114.8000 142.2000 115.6000 145.0000 ;
	    RECT 116.4000 142.2000 117.2000 145.0000 ;
	    RECT 118.0000 142.2000 118.8000 145.0000 ;
	    RECT 119.6000 142.2000 120.4000 145.0000 ;
	    RECT 121.2000 142.2000 122.0000 145.4000 ;
	    RECT 127.6000 142.2000 128.4000 147.4000 ;
	    RECT 129.4000 146.8000 130.2000 151.2000 ;
	    RECT 134.4000 148.4000 135.0000 151.8000 ;
	    RECT 135.6000 148.8000 136.4000 150.4000 ;
	    RECT 130.8000 148.3000 131.6000 148.4000 ;
	    RECT 132.4000 148.3000 135.0000 148.4000 ;
	    RECT 130.8000 147.7000 135.0000 148.3000 ;
	    RECT 137.2000 148.3000 138.0000 148.4000 ;
	    RECT 138.8000 148.3000 139.6000 159.8000 ;
	    RECT 140.4000 152.3000 141.2000 152.4000 ;
	    RECT 142.0000 152.3000 142.8000 159.8000 ;
	    RECT 146.8000 155.8000 147.6000 159.8000 ;
	    RECT 140.4000 151.7000 142.8000 152.3000 ;
	    RECT 140.4000 151.6000 141.2000 151.7000 ;
	    RECT 137.2000 148.2000 139.6000 148.3000 ;
	    RECT 130.8000 147.6000 131.6000 147.7000 ;
	    RECT 132.4000 147.6000 135.0000 147.7000 ;
	    RECT 136.4000 147.7000 139.6000 148.2000 ;
	    RECT 136.4000 147.6000 138.0000 147.7000 ;
	    RECT 129.2000 146.0000 130.2000 146.8000 ;
	    RECT 132.6000 146.2000 133.2000 147.6000 ;
	    RECT 136.4000 147.2000 137.2000 147.6000 ;
	    RECT 134.2000 146.2000 137.8000 146.6000 ;
	    RECT 129.2000 142.2000 130.0000 146.0000 ;
	    RECT 132.4000 142.2000 133.2000 146.2000 ;
	    RECT 134.0000 146.0000 138.0000 146.2000 ;
	    RECT 134.0000 142.2000 134.8000 146.0000 ;
	    RECT 137.2000 142.2000 138.0000 146.0000 ;
	    RECT 138.8000 142.2000 139.6000 147.7000 ;
	    RECT 140.4000 144.8000 141.2000 146.4000 ;
	    RECT 142.0000 142.2000 142.8000 151.7000 ;
	    RECT 147.0000 151.6000 147.6000 155.8000 ;
	    RECT 150.0000 151.8000 150.8000 159.8000 ;
	    RECT 151.6000 152.4000 152.4000 159.8000 ;
	    RECT 154.8000 158.3000 155.6000 159.8000 ;
	    RECT 159.6000 158.3000 160.4000 158.4000 ;
	    RECT 154.8000 157.7000 160.4000 158.3000 ;
	    RECT 151.6000 151.8000 153.8000 152.4000 ;
	    RECT 154.8000 151.8000 155.6000 157.7000 ;
	    RECT 159.6000 157.6000 160.4000 157.7000 ;
	    RECT 147.0000 151.0000 149.4000 151.6000 ;
	    RECT 146.8000 149.6000 147.6000 150.4000 ;
	    RECT 145.2000 147.6000 146.0000 149.2000 ;
	    RECT 147.0000 148.8000 147.6000 149.6000 ;
	    RECT 147.0000 148.2000 148.0000 148.8000 ;
	    RECT 147.2000 148.0000 148.0000 148.2000 ;
	    RECT 148.8000 147.6000 149.4000 151.0000 ;
	    RECT 150.2000 150.4000 150.8000 151.8000 ;
	    RECT 153.2000 151.2000 153.8000 151.8000 ;
	    RECT 153.2000 150.4000 154.4000 151.2000 ;
	    RECT 150.0000 149.6000 150.8000 150.4000 ;
	    RECT 148.8000 147.4000 149.6000 147.6000 ;
	    RECT 146.6000 147.0000 149.6000 147.4000 ;
	    RECT 145.4000 146.8000 149.6000 147.0000 ;
	    RECT 145.4000 146.4000 147.2000 146.8000 ;
	    RECT 143.6000 144.8000 144.4000 146.4000 ;
	    RECT 145.4000 146.2000 146.0000 146.4000 ;
	    RECT 150.2000 146.2000 150.8000 149.6000 ;
	    RECT 151.6000 148.8000 152.4000 150.4000 ;
	    RECT 153.2000 147.4000 153.8000 150.4000 ;
	    RECT 155.0000 149.6000 155.6000 151.8000 ;
	    RECT 162.8000 151.2000 163.6000 159.8000 ;
	    RECT 166.0000 151.2000 166.8000 159.8000 ;
	    RECT 169.2000 151.2000 170.0000 159.8000 ;
	    RECT 172.4000 151.2000 173.2000 159.8000 ;
	    RECT 175.6000 152.4000 176.4000 159.8000 ;
	    RECT 178.8000 152.4000 179.6000 159.8000 ;
	    RECT 175.6000 151.8000 179.6000 152.4000 ;
	    RECT 180.4000 151.8000 181.2000 159.8000 ;
	    RECT 162.8000 150.4000 164.6000 151.2000 ;
	    RECT 166.0000 150.4000 168.2000 151.2000 ;
	    RECT 169.2000 150.4000 171.4000 151.2000 ;
	    RECT 172.4000 150.4000 174.8000 151.2000 ;
	    RECT 176.4000 150.4000 177.2000 150.8000 ;
	    RECT 180.4000 150.4000 181.0000 151.8000 ;
	    RECT 145.2000 142.2000 146.0000 146.2000 ;
	    RECT 149.4000 145.2000 150.8000 146.2000 ;
	    RECT 151.6000 146.8000 153.8000 147.4000 ;
	    RECT 149.4000 144.4000 150.2000 145.2000 ;
	    RECT 149.4000 143.6000 150.8000 144.4000 ;
	    RECT 149.4000 142.2000 150.2000 143.6000 ;
	    RECT 151.6000 142.2000 152.4000 146.8000 ;
	    RECT 154.8000 142.2000 155.6000 149.6000 ;
	    RECT 163.8000 149.0000 164.6000 150.4000 ;
	    RECT 167.4000 149.0000 168.2000 150.4000 ;
	    RECT 170.6000 149.0000 171.4000 150.4000 ;
	    RECT 163.8000 148.2000 166.4000 149.0000 ;
	    RECT 167.4000 148.2000 169.8000 149.0000 ;
	    RECT 170.6000 148.2000 173.2000 149.0000 ;
	    RECT 163.8000 147.6000 164.6000 148.2000 ;
	    RECT 167.4000 147.6000 168.2000 148.2000 ;
	    RECT 170.6000 147.6000 171.4000 148.2000 ;
	    RECT 174.0000 147.6000 174.8000 150.4000 ;
	    RECT 175.6000 149.8000 177.2000 150.4000 ;
	    RECT 178.8000 149.8000 181.2000 150.4000 ;
	    RECT 175.6000 149.6000 176.4000 149.8000 ;
	    RECT 177.2000 147.6000 178.0000 149.2000 ;
	    RECT 162.8000 146.8000 164.6000 147.6000 ;
	    RECT 166.0000 146.8000 168.2000 147.6000 ;
	    RECT 169.2000 146.8000 171.4000 147.6000 ;
	    RECT 172.4000 146.8000 174.8000 147.6000 ;
	    RECT 162.8000 142.2000 163.6000 146.8000 ;
	    RECT 166.0000 142.2000 166.8000 146.8000 ;
	    RECT 169.2000 142.2000 170.0000 146.8000 ;
	    RECT 172.4000 142.2000 173.2000 146.8000 ;
	    RECT 178.8000 146.2000 179.4000 149.8000 ;
	    RECT 180.4000 149.6000 181.2000 149.8000 ;
	    RECT 180.4000 148.3000 181.2000 148.4000 ;
	    RECT 182.0000 148.3000 182.8000 159.8000 ;
	    RECT 186.8000 156.4000 187.6000 159.8000 ;
	    RECT 186.6000 155.8000 187.6000 156.4000 ;
	    RECT 186.6000 155.2000 187.2000 155.8000 ;
	    RECT 190.0000 155.2000 190.8000 159.8000 ;
	    RECT 193.2000 157.0000 194.0000 159.8000 ;
	    RECT 194.8000 157.0000 195.6000 159.8000 ;
	    RECT 180.4000 147.7000 182.8000 148.3000 ;
	    RECT 180.4000 147.6000 181.2000 147.7000 ;
	    RECT 178.8000 142.2000 179.6000 146.2000 ;
	    RECT 180.4000 145.6000 181.2000 146.4000 ;
	    RECT 180.2000 144.8000 181.0000 145.6000 ;
	    RECT 182.0000 142.2000 182.8000 147.7000 ;
	    RECT 185.2000 154.6000 187.2000 155.2000 ;
	    RECT 185.2000 149.0000 186.0000 154.6000 ;
	    RECT 187.8000 154.4000 192.0000 155.2000 ;
	    RECT 196.4000 155.0000 197.2000 159.8000 ;
	    RECT 199.6000 155.0000 200.4000 159.8000 ;
	    RECT 187.8000 154.0000 188.4000 154.4000 ;
	    RECT 186.8000 153.2000 188.4000 154.0000 ;
	    RECT 191.4000 153.8000 197.2000 154.4000 ;
	    RECT 189.4000 153.2000 190.8000 153.8000 ;
	    RECT 189.4000 153.0000 195.6000 153.2000 ;
	    RECT 190.2000 152.6000 195.6000 153.0000 ;
	    RECT 194.8000 152.4000 195.6000 152.6000 ;
	    RECT 196.6000 153.0000 197.2000 153.8000 ;
	    RECT 197.8000 153.6000 200.4000 154.4000 ;
	    RECT 202.8000 153.6000 203.6000 159.8000 ;
	    RECT 204.4000 157.0000 205.2000 159.8000 ;
	    RECT 206.0000 157.0000 206.8000 159.8000 ;
	    RECT 207.6000 157.0000 208.4000 159.8000 ;
	    RECT 206.0000 154.4000 210.2000 155.2000 ;
	    RECT 210.8000 154.4000 211.6000 159.8000 ;
	    RECT 214.0000 155.2000 214.8000 159.8000 ;
	    RECT 214.0000 154.6000 216.6000 155.2000 ;
	    RECT 210.8000 153.6000 213.4000 154.4000 ;
	    RECT 204.4000 153.0000 205.2000 153.2000 ;
	    RECT 196.6000 152.4000 205.2000 153.0000 ;
	    RECT 207.6000 153.0000 208.4000 153.2000 ;
	    RECT 216.0000 153.0000 216.6000 154.6000 ;
	    RECT 207.6000 152.4000 216.6000 153.0000 ;
	    RECT 216.0000 150.6000 216.6000 152.4000 ;
	    RECT 217.2000 152.0000 218.0000 159.8000 ;
	    RECT 220.4000 152.4000 221.2000 159.8000 ;
	    RECT 217.2000 151.2000 218.2000 152.0000 ;
	    RECT 220.4000 151.8000 222.6000 152.4000 ;
	    RECT 186.6000 150.0000 210.0000 150.6000 ;
	    RECT 216.0000 150.0000 216.8000 150.6000 ;
	    RECT 186.6000 149.8000 187.4000 150.0000 ;
	    RECT 188.4000 149.6000 189.2000 150.0000 ;
	    RECT 190.0000 149.6000 190.8000 150.0000 ;
	    RECT 191.6000 149.6000 192.4000 150.0000 ;
	    RECT 209.2000 149.4000 210.0000 150.0000 ;
	    RECT 185.2000 148.2000 194.0000 149.0000 ;
	    RECT 194.6000 148.6000 196.6000 149.4000 ;
	    RECT 200.4000 148.6000 203.6000 149.4000 ;
	    RECT 183.6000 144.8000 184.4000 146.4000 ;
	    RECT 185.2000 142.2000 186.0000 148.2000 ;
	    RECT 187.6000 146.8000 190.6000 147.6000 ;
	    RECT 189.8000 146.2000 190.6000 146.8000 ;
	    RECT 195.8000 146.2000 196.6000 148.6000 ;
	    RECT 198.0000 146.8000 198.8000 148.4000 ;
	    RECT 203.2000 147.8000 204.0000 148.0000 ;
	    RECT 199.6000 147.2000 204.0000 147.8000 ;
	    RECT 199.6000 147.0000 200.4000 147.2000 ;
	    RECT 206.0000 146.4000 206.8000 149.2000 ;
	    RECT 211.8000 148.6000 215.6000 149.4000 ;
	    RECT 211.8000 147.4000 212.6000 148.6000 ;
	    RECT 216.2000 148.0000 216.8000 150.0000 ;
	    RECT 199.6000 146.2000 200.4000 146.4000 ;
	    RECT 189.8000 145.4000 192.4000 146.2000 ;
	    RECT 195.8000 145.6000 200.4000 146.2000 ;
	    RECT 201.2000 145.6000 202.8000 146.4000 ;
	    RECT 205.8000 145.6000 206.8000 146.4000 ;
	    RECT 210.8000 146.8000 212.6000 147.4000 ;
	    RECT 215.6000 147.4000 216.8000 148.0000 ;
	    RECT 217.4000 150.3000 218.2000 151.2000 ;
	    RECT 222.0000 151.2000 222.6000 151.8000 ;
	    RECT 222.0000 150.4000 223.2000 151.2000 ;
	    RECT 220.4000 150.3000 221.2000 150.4000 ;
	    RECT 217.4000 149.7000 221.2000 150.3000 ;
	    RECT 210.8000 146.2000 211.6000 146.8000 ;
	    RECT 191.6000 142.2000 192.4000 145.4000 ;
	    RECT 209.2000 145.4000 211.6000 146.2000 ;
	    RECT 193.2000 142.2000 194.0000 145.0000 ;
	    RECT 194.8000 142.2000 195.6000 145.0000 ;
	    RECT 196.4000 142.2000 197.2000 145.0000 ;
	    RECT 199.6000 142.2000 200.4000 145.0000 ;
	    RECT 202.8000 142.2000 203.6000 145.0000 ;
	    RECT 204.4000 142.2000 205.2000 145.0000 ;
	    RECT 206.0000 142.2000 206.8000 145.0000 ;
	    RECT 207.6000 142.2000 208.4000 145.0000 ;
	    RECT 209.2000 142.2000 210.0000 145.4000 ;
	    RECT 215.6000 142.2000 216.4000 147.4000 ;
	    RECT 217.4000 146.8000 218.2000 149.7000 ;
	    RECT 220.4000 148.8000 221.2000 149.7000 ;
	    RECT 222.0000 147.4000 222.6000 150.4000 ;
	    RECT 217.2000 146.0000 218.2000 146.8000 ;
	    RECT 220.4000 146.8000 222.6000 147.4000 ;
	    RECT 217.2000 142.2000 218.0000 146.0000 ;
	    RECT 220.4000 142.2000 221.2000 146.8000 ;
	    RECT 4.4000 135.2000 5.2000 139.8000 ;
	    RECT 6.0000 135.6000 6.8000 137.2000 ;
	    RECT 3.0000 134.6000 5.2000 135.2000 ;
	    RECT 3.0000 131.6000 3.6000 134.6000 ;
	    RECT 4.4000 131.6000 5.2000 133.2000 ;
	    RECT 7.6000 132.3000 8.4000 139.8000 ;
	    RECT 13.0000 138.4000 13.8000 139.0000 ;
	    RECT 13.0000 137.6000 14.8000 138.4000 ;
	    RECT 13.0000 136.0000 13.8000 137.6000 ;
	    RECT 17.2000 137.0000 18.0000 139.0000 ;
	    RECT 12.2000 135.4000 13.8000 136.0000 ;
	    RECT 12.2000 135.0000 13.0000 135.4000 ;
	    RECT 12.2000 134.4000 12.8000 135.0000 ;
	    RECT 17.4000 134.8000 18.0000 137.0000 ;
	    RECT 20.4000 136.0000 21.2000 139.8000 ;
	    RECT 10.8000 133.6000 12.8000 134.4000 ;
	    RECT 13.8000 134.2000 18.0000 134.8000 ;
	    RECT 20.2000 135.2000 21.2000 136.0000 ;
	    RECT 13.8000 133.8000 14.8000 134.2000 ;
	    RECT 10.8000 132.3000 11.6000 132.4000 ;
	    RECT 7.6000 131.7000 11.6000 132.3000 ;
	    RECT 2.4000 130.8000 3.6000 131.6000 ;
	    RECT 3.0000 130.2000 3.6000 130.8000 ;
	    RECT 3.0000 129.6000 5.2000 130.2000 ;
	    RECT 4.4000 122.2000 5.2000 129.6000 ;
	    RECT 7.6000 122.2000 8.4000 131.7000 ;
	    RECT 10.8000 130.8000 11.6000 131.7000 ;
	    RECT 12.2000 129.8000 12.8000 133.6000 ;
	    RECT 13.4000 133.0000 14.8000 133.8000 ;
	    RECT 14.2000 131.0000 14.8000 133.0000 ;
	    RECT 15.6000 131.6000 16.4000 133.2000 ;
	    RECT 17.2000 131.6000 18.0000 133.2000 ;
	    RECT 14.2000 130.4000 18.0000 131.0000 ;
	    RECT 12.2000 129.2000 13.8000 129.8000 ;
	    RECT 13.0000 122.2000 13.8000 129.2000 ;
	    RECT 17.4000 127.0000 18.0000 130.4000 ;
	    RECT 20.2000 130.8000 21.0000 135.2000 ;
	    RECT 22.0000 134.6000 22.8000 139.8000 ;
	    RECT 28.4000 136.6000 29.2000 139.8000 ;
	    RECT 30.0000 137.0000 30.8000 139.8000 ;
	    RECT 31.6000 137.0000 32.4000 139.8000 ;
	    RECT 33.2000 137.0000 34.0000 139.8000 ;
	    RECT 34.8000 137.0000 35.6000 139.8000 ;
	    RECT 38.0000 137.0000 38.8000 139.8000 ;
	    RECT 41.2000 137.0000 42.0000 139.8000 ;
	    RECT 42.8000 137.0000 43.6000 139.8000 ;
	    RECT 44.4000 137.0000 45.2000 139.8000 ;
	    RECT 26.8000 135.8000 29.2000 136.6000 ;
	    RECT 46.0000 136.6000 46.8000 139.8000 ;
	    RECT 26.8000 135.2000 27.6000 135.8000 ;
	    RECT 21.6000 134.0000 22.8000 134.6000 ;
	    RECT 25.8000 134.6000 27.6000 135.2000 ;
	    RECT 31.6000 135.6000 32.6000 136.4000 ;
	    RECT 35.6000 135.6000 37.2000 136.4000 ;
	    RECT 38.0000 135.8000 42.6000 136.4000 ;
	    RECT 46.0000 135.8000 48.6000 136.6000 ;
	    RECT 38.0000 135.6000 38.8000 135.8000 ;
	    RECT 21.6000 132.0000 22.2000 134.0000 ;
	    RECT 25.8000 133.4000 26.6000 134.6000 ;
	    RECT 22.8000 132.6000 26.6000 133.4000 ;
	    RECT 31.6000 132.8000 32.4000 135.6000 ;
	    RECT 38.0000 134.8000 38.8000 135.0000 ;
	    RECT 34.4000 134.2000 38.8000 134.8000 ;
	    RECT 34.4000 134.0000 35.2000 134.2000 ;
	    RECT 39.6000 133.6000 40.4000 135.2000 ;
	    RECT 41.8000 133.4000 42.6000 135.8000 ;
	    RECT 47.8000 135.2000 48.6000 135.8000 ;
	    RECT 47.8000 134.4000 50.8000 135.2000 ;
	    RECT 52.4000 133.8000 53.2000 139.8000 ;
	    RECT 54.0000 136.0000 54.8000 139.8000 ;
	    RECT 57.2000 136.0000 58.0000 139.8000 ;
	    RECT 54.0000 135.8000 58.0000 136.0000 ;
	    RECT 54.2000 135.4000 57.8000 135.8000 ;
	    RECT 58.8000 135.6000 59.6000 139.8000 ;
	    RECT 54.8000 134.4000 55.6000 134.8000 ;
	    RECT 58.8000 134.4000 59.4000 135.6000 ;
	    RECT 34.8000 132.6000 38.0000 133.4000 ;
	    RECT 41.8000 132.6000 43.8000 133.4000 ;
	    RECT 44.4000 133.0000 53.2000 133.8000 ;
	    RECT 54.0000 133.8000 55.6000 134.4000 ;
	    RECT 54.0000 133.6000 54.8000 133.8000 ;
	    RECT 57.0000 133.6000 59.6000 134.4000 ;
	    RECT 28.4000 132.0000 29.2000 132.6000 ;
	    RECT 46.0000 132.0000 46.8000 132.4000 ;
	    RECT 51.0000 132.0000 51.8000 132.2000 ;
	    RECT 21.6000 131.4000 22.4000 132.0000 ;
	    RECT 28.4000 131.4000 51.8000 132.0000 ;
	    RECT 20.2000 130.0000 21.2000 130.8000 ;
	    RECT 17.2000 123.0000 18.0000 127.0000 ;
	    RECT 20.4000 122.2000 21.2000 130.0000 ;
	    RECT 21.8000 129.6000 22.4000 131.4000 ;
	    RECT 21.8000 129.0000 30.8000 129.6000 ;
	    RECT 21.8000 127.4000 22.4000 129.0000 ;
	    RECT 30.0000 128.8000 30.8000 129.0000 ;
	    RECT 33.2000 129.0000 41.8000 129.6000 ;
	    RECT 33.2000 128.8000 34.0000 129.0000 ;
	    RECT 25.0000 127.6000 27.6000 128.4000 ;
	    RECT 21.8000 126.8000 24.4000 127.4000 ;
	    RECT 23.6000 122.2000 24.4000 126.8000 ;
	    RECT 26.8000 122.2000 27.6000 127.6000 ;
	    RECT 28.2000 126.8000 32.4000 127.6000 ;
	    RECT 30.0000 122.2000 30.8000 125.0000 ;
	    RECT 31.6000 122.2000 32.4000 125.0000 ;
	    RECT 33.2000 122.2000 34.0000 125.0000 ;
	    RECT 34.8000 122.2000 35.6000 128.4000 ;
	    RECT 38.0000 127.6000 40.6000 128.4000 ;
	    RECT 41.2000 128.2000 41.8000 129.0000 ;
	    RECT 42.8000 129.4000 43.6000 129.6000 ;
	    RECT 42.8000 129.0000 48.2000 129.4000 ;
	    RECT 42.8000 128.8000 49.0000 129.0000 ;
	    RECT 47.6000 128.2000 49.0000 128.8000 ;
	    RECT 41.2000 127.6000 47.0000 128.2000 ;
	    RECT 50.0000 128.0000 51.6000 128.8000 ;
	    RECT 50.0000 127.6000 50.6000 128.0000 ;
	    RECT 38.0000 122.2000 38.8000 127.0000 ;
	    RECT 41.2000 122.2000 42.0000 127.0000 ;
	    RECT 46.4000 126.8000 50.6000 127.6000 ;
	    RECT 52.4000 127.4000 53.2000 133.0000 ;
	    RECT 55.6000 131.6000 56.4000 133.2000 ;
	    RECT 57.0000 130.2000 57.6000 133.6000 ;
	    RECT 60.4000 132.4000 61.2000 139.8000 ;
	    RECT 63.6000 135.2000 64.4000 139.8000 ;
	    RECT 62.2000 134.6000 64.4000 135.2000 ;
	    RECT 70.0000 135.2000 70.8000 139.8000 ;
	    RECT 70.0000 134.6000 72.2000 135.2000 ;
	    RECT 58.8000 130.2000 59.6000 130.4000 ;
	    RECT 51.2000 126.8000 53.2000 127.4000 ;
	    RECT 56.6000 129.6000 57.6000 130.2000 ;
	    RECT 58.2000 129.6000 59.6000 130.2000 ;
	    RECT 60.4000 130.2000 61.0000 132.4000 ;
	    RECT 62.2000 131.6000 62.8000 134.6000 ;
	    RECT 63.6000 132.3000 64.4000 133.2000 ;
	    RECT 70.0000 132.3000 70.8000 133.2000 ;
	    RECT 63.6000 131.7000 70.8000 132.3000 ;
	    RECT 63.6000 131.6000 64.4000 131.7000 ;
	    RECT 70.0000 131.6000 70.8000 131.7000 ;
	    RECT 71.6000 131.6000 72.2000 134.6000 ;
	    RECT 73.2000 134.3000 74.0000 139.8000 ;
	    RECT 75.0000 136.4000 75.8000 137.2000 ;
	    RECT 74.8000 135.6000 75.6000 136.4000 ;
	    RECT 76.4000 135.8000 77.2000 139.8000 ;
	    RECT 74.8000 134.3000 75.6000 134.4000 ;
	    RECT 73.2000 133.7000 75.6000 134.3000 ;
	    RECT 73.2000 132.4000 74.0000 133.7000 ;
	    RECT 74.8000 133.6000 75.6000 133.7000 ;
	    RECT 61.6000 130.8000 62.8000 131.6000 ;
	    RECT 62.2000 130.2000 62.8000 130.8000 ;
	    RECT 71.6000 130.8000 72.8000 131.6000 ;
	    RECT 71.6000 130.2000 72.2000 130.8000 ;
	    RECT 73.4000 130.2000 74.0000 132.4000 ;
	    RECT 74.8000 132.2000 75.6000 132.4000 ;
	    RECT 76.6000 132.2000 77.2000 135.8000 ;
	    RECT 81.2000 137.0000 82.0000 139.0000 ;
	    RECT 85.4000 138.4000 86.2000 139.0000 ;
	    RECT 84.4000 137.6000 86.2000 138.4000 ;
	    RECT 81.2000 134.8000 81.8000 137.0000 ;
	    RECT 85.4000 136.0000 86.2000 137.6000 ;
	    RECT 85.4000 135.4000 87.0000 136.0000 ;
	    RECT 86.2000 135.0000 87.0000 135.4000 ;
	    RECT 78.0000 132.8000 78.8000 134.4000 ;
	    RECT 81.2000 134.2000 85.4000 134.8000 ;
	    RECT 84.4000 133.8000 85.4000 134.2000 ;
	    RECT 86.4000 134.4000 87.0000 135.0000 ;
	    RECT 79.6000 132.2000 80.4000 132.4000 ;
	    RECT 74.8000 131.6000 77.2000 132.2000 ;
	    RECT 78.8000 131.6000 80.4000 132.2000 ;
	    RECT 81.2000 131.6000 82.0000 133.2000 ;
	    RECT 82.8000 131.6000 83.6000 133.2000 ;
	    RECT 84.4000 133.0000 85.8000 133.8000 ;
	    RECT 86.4000 133.6000 88.4000 134.4000 ;
	    RECT 75.0000 130.2000 75.6000 131.6000 ;
	    RECT 78.8000 131.2000 79.6000 131.6000 ;
	    RECT 84.4000 131.0000 85.0000 133.0000 ;
	    RECT 81.2000 130.4000 85.0000 131.0000 ;
	    RECT 42.8000 122.2000 43.6000 125.0000 ;
	    RECT 44.4000 122.2000 45.2000 125.0000 ;
	    RECT 47.6000 122.2000 48.4000 126.8000 ;
	    RECT 51.2000 126.2000 51.8000 126.8000 ;
	    RECT 50.8000 125.6000 51.8000 126.2000 ;
	    RECT 50.8000 122.2000 51.6000 125.6000 ;
	    RECT 56.6000 122.2000 57.4000 129.6000 ;
	    RECT 58.2000 128.4000 58.8000 129.6000 ;
	    RECT 58.0000 127.6000 58.8000 128.4000 ;
	    RECT 60.4000 122.2000 61.2000 130.2000 ;
	    RECT 62.2000 129.6000 64.4000 130.2000 ;
	    RECT 63.6000 122.2000 64.4000 129.6000 ;
	    RECT 70.0000 129.6000 72.2000 130.2000 ;
	    RECT 70.0000 122.2000 70.8000 129.6000 ;
	    RECT 73.2000 122.2000 74.0000 130.2000 ;
	    RECT 74.8000 122.2000 75.6000 130.2000 ;
	    RECT 76.4000 129.6000 80.4000 130.2000 ;
	    RECT 76.4000 122.2000 77.2000 129.6000 ;
	    RECT 79.6000 122.2000 80.4000 129.6000 ;
	    RECT 81.2000 127.0000 81.8000 130.4000 ;
	    RECT 86.4000 129.8000 87.0000 133.6000 ;
	    RECT 87.6000 132.3000 88.4000 132.4000 ;
	    RECT 90.8000 132.3000 91.6000 139.8000 ;
	    RECT 92.4000 135.6000 93.2000 137.2000 ;
	    RECT 95.6000 135.2000 96.4000 139.8000 ;
	    RECT 98.8000 135.2000 99.6000 139.8000 ;
	    RECT 102.0000 135.2000 102.8000 139.8000 ;
	    RECT 105.2000 135.2000 106.0000 139.8000 ;
	    RECT 87.6000 131.7000 91.6000 132.3000 ;
	    RECT 87.6000 130.8000 88.4000 131.7000 ;
	    RECT 85.4000 129.2000 87.0000 129.8000 ;
	    RECT 81.2000 123.0000 82.0000 127.0000 ;
	    RECT 85.4000 122.2000 86.2000 129.2000 ;
	    RECT 90.8000 122.2000 91.6000 131.7000 ;
	    RECT 94.0000 134.4000 96.4000 135.2000 ;
	    RECT 97.4000 134.4000 99.6000 135.2000 ;
	    RECT 100.6000 134.4000 102.8000 135.2000 ;
	    RECT 104.2000 134.4000 106.0000 135.2000 ;
	    RECT 94.0000 131.6000 94.8000 134.4000 ;
	    RECT 97.4000 133.8000 98.2000 134.4000 ;
	    RECT 100.6000 133.8000 101.4000 134.4000 ;
	    RECT 104.2000 133.8000 105.0000 134.4000 ;
	    RECT 95.6000 133.0000 98.2000 133.8000 ;
	    RECT 99.0000 133.0000 101.4000 133.8000 ;
	    RECT 102.4000 133.0000 105.0000 133.8000 ;
	    RECT 97.4000 131.6000 98.2000 133.0000 ;
	    RECT 100.6000 131.6000 101.4000 133.0000 ;
	    RECT 104.2000 131.6000 105.0000 133.0000 ;
	    RECT 108.4000 133.8000 109.2000 139.8000 ;
	    RECT 114.8000 136.6000 115.6000 139.8000 ;
	    RECT 116.4000 137.0000 117.2000 139.8000 ;
	    RECT 118.0000 137.0000 118.8000 139.8000 ;
	    RECT 119.6000 137.0000 120.4000 139.8000 ;
	    RECT 122.8000 137.0000 123.6000 139.8000 ;
	    RECT 126.0000 137.0000 126.8000 139.8000 ;
	    RECT 127.6000 137.0000 128.4000 139.8000 ;
	    RECT 129.2000 137.0000 130.0000 139.8000 ;
	    RECT 130.8000 137.0000 131.6000 139.8000 ;
	    RECT 113.0000 135.8000 115.6000 136.6000 ;
	    RECT 132.4000 136.6000 133.2000 139.8000 ;
	    RECT 119.0000 135.8000 123.6000 136.4000 ;
	    RECT 113.0000 135.2000 113.8000 135.8000 ;
	    RECT 110.8000 134.4000 113.8000 135.2000 ;
	    RECT 108.4000 133.0000 117.2000 133.8000 ;
	    RECT 119.0000 133.4000 119.8000 135.8000 ;
	    RECT 122.8000 135.6000 123.6000 135.8000 ;
	    RECT 124.4000 135.6000 126.0000 136.4000 ;
	    RECT 129.0000 135.6000 130.0000 136.4000 ;
	    RECT 132.4000 135.8000 134.8000 136.6000 ;
	    RECT 121.2000 133.6000 122.0000 135.2000 ;
	    RECT 122.8000 134.8000 123.6000 135.0000 ;
	    RECT 122.8000 134.2000 127.2000 134.8000 ;
	    RECT 126.4000 134.0000 127.2000 134.2000 ;
	    RECT 94.0000 130.8000 96.4000 131.6000 ;
	    RECT 97.4000 130.8000 99.6000 131.6000 ;
	    RECT 100.6000 130.8000 102.8000 131.6000 ;
	    RECT 104.2000 130.8000 106.0000 131.6000 ;
	    RECT 95.6000 122.2000 96.4000 130.8000 ;
	    RECT 98.8000 122.2000 99.6000 130.8000 ;
	    RECT 102.0000 122.2000 102.8000 130.8000 ;
	    RECT 105.2000 122.2000 106.0000 130.8000 ;
	    RECT 108.4000 127.4000 109.2000 133.0000 ;
	    RECT 117.8000 132.6000 119.8000 133.4000 ;
	    RECT 123.6000 132.6000 126.8000 133.4000 ;
	    RECT 129.2000 132.8000 130.0000 135.6000 ;
	    RECT 134.0000 135.2000 134.8000 135.8000 ;
	    RECT 134.0000 134.6000 135.8000 135.2000 ;
	    RECT 135.0000 133.4000 135.8000 134.6000 ;
	    RECT 138.8000 134.6000 139.6000 139.8000 ;
	    RECT 140.4000 136.3000 141.2000 139.8000 ;
	    RECT 145.2000 138.3000 146.0000 139.8000 ;
	    RECT 146.8000 138.3000 147.6000 138.4000 ;
	    RECT 145.2000 137.7000 147.6000 138.3000 ;
	    RECT 142.0000 136.3000 142.8000 136.4000 ;
	    RECT 140.4000 135.7000 142.8000 136.3000 ;
	    RECT 140.4000 135.2000 141.4000 135.7000 ;
	    RECT 142.0000 135.6000 142.8000 135.7000 ;
	    RECT 143.6000 135.6000 144.4000 137.2000 ;
	    RECT 138.8000 134.0000 140.0000 134.6000 ;
	    RECT 135.0000 132.6000 138.8000 133.4000 ;
	    RECT 109.8000 132.0000 110.6000 132.2000 ;
	    RECT 111.6000 132.0000 112.4000 132.4000 ;
	    RECT 114.8000 132.0000 115.6000 132.4000 ;
	    RECT 132.4000 132.0000 133.2000 132.6000 ;
	    RECT 139.4000 132.0000 140.0000 134.0000 ;
	    RECT 109.8000 131.4000 133.2000 132.0000 ;
	    RECT 139.2000 131.4000 140.0000 132.0000 ;
	    RECT 139.2000 129.6000 139.8000 131.4000 ;
	    RECT 140.6000 130.8000 141.4000 135.2000 ;
	    RECT 118.0000 129.4000 118.8000 129.6000 ;
	    RECT 113.4000 129.0000 118.8000 129.4000 ;
	    RECT 112.6000 128.8000 118.8000 129.0000 ;
	    RECT 119.8000 129.0000 128.4000 129.6000 ;
	    RECT 110.0000 128.0000 111.6000 128.8000 ;
	    RECT 112.6000 128.2000 114.0000 128.8000 ;
	    RECT 119.8000 128.2000 120.4000 129.0000 ;
	    RECT 127.6000 128.8000 128.4000 129.0000 ;
	    RECT 130.8000 129.0000 139.8000 129.6000 ;
	    RECT 130.8000 128.8000 131.6000 129.0000 ;
	    RECT 111.0000 127.6000 111.6000 128.0000 ;
	    RECT 114.6000 127.6000 120.4000 128.2000 ;
	    RECT 121.0000 127.6000 123.6000 128.4000 ;
	    RECT 108.4000 126.8000 110.4000 127.4000 ;
	    RECT 111.0000 126.8000 115.2000 127.6000 ;
	    RECT 109.8000 126.2000 110.4000 126.8000 ;
	    RECT 109.8000 125.6000 110.8000 126.2000 ;
	    RECT 110.0000 122.2000 110.8000 125.6000 ;
	    RECT 113.2000 122.2000 114.0000 126.8000 ;
	    RECT 116.4000 122.2000 117.2000 125.0000 ;
	    RECT 118.0000 122.2000 118.8000 125.0000 ;
	    RECT 119.6000 122.2000 120.4000 127.0000 ;
	    RECT 122.8000 122.2000 123.6000 127.0000 ;
	    RECT 126.0000 122.2000 126.8000 128.4000 ;
	    RECT 134.0000 127.6000 136.6000 128.4000 ;
	    RECT 129.2000 126.8000 133.4000 127.6000 ;
	    RECT 127.6000 122.2000 128.4000 125.0000 ;
	    RECT 129.2000 122.2000 130.0000 125.0000 ;
	    RECT 130.8000 122.2000 131.6000 125.0000 ;
	    RECT 134.0000 122.2000 134.8000 127.6000 ;
	    RECT 139.2000 127.4000 139.8000 129.0000 ;
	    RECT 137.2000 126.8000 139.8000 127.4000 ;
	    RECT 140.4000 130.0000 141.4000 130.8000 ;
	    RECT 137.2000 122.2000 138.0000 126.8000 ;
	    RECT 140.4000 122.2000 141.2000 130.0000 ;
	    RECT 145.2000 122.2000 146.0000 137.7000 ;
	    RECT 146.8000 137.6000 147.6000 137.7000 ;
	    RECT 151.6000 133.8000 152.4000 139.8000 ;
	    RECT 158.0000 136.6000 158.8000 139.8000 ;
	    RECT 159.6000 137.0000 160.4000 139.8000 ;
	    RECT 161.2000 137.0000 162.0000 139.8000 ;
	    RECT 162.8000 137.0000 163.6000 139.8000 ;
	    RECT 166.0000 137.0000 166.8000 139.8000 ;
	    RECT 169.2000 137.0000 170.0000 139.8000 ;
	    RECT 170.8000 137.0000 171.6000 139.8000 ;
	    RECT 172.4000 137.0000 173.2000 139.8000 ;
	    RECT 174.0000 137.0000 174.8000 139.8000 ;
	    RECT 156.2000 135.8000 158.8000 136.6000 ;
	    RECT 175.6000 136.6000 176.4000 139.8000 ;
	    RECT 162.2000 135.8000 166.8000 136.4000 ;
	    RECT 156.2000 135.2000 157.0000 135.8000 ;
	    RECT 154.0000 134.4000 157.0000 135.2000 ;
	    RECT 151.6000 133.0000 160.4000 133.8000 ;
	    RECT 162.2000 133.4000 163.0000 135.8000 ;
	    RECT 166.0000 135.6000 166.8000 135.8000 ;
	    RECT 167.6000 135.6000 169.2000 136.4000 ;
	    RECT 172.2000 135.6000 173.2000 136.4000 ;
	    RECT 175.6000 135.8000 178.0000 136.6000 ;
	    RECT 164.4000 133.6000 165.2000 135.2000 ;
	    RECT 166.0000 134.8000 166.8000 135.0000 ;
	    RECT 166.0000 134.2000 170.4000 134.8000 ;
	    RECT 169.6000 134.0000 170.4000 134.2000 ;
	    RECT 151.6000 127.4000 152.4000 133.0000 ;
	    RECT 161.0000 132.6000 163.0000 133.4000 ;
	    RECT 166.8000 132.6000 170.0000 133.4000 ;
	    RECT 172.4000 132.8000 173.2000 135.6000 ;
	    RECT 177.2000 135.2000 178.0000 135.8000 ;
	    RECT 177.2000 134.6000 179.0000 135.2000 ;
	    RECT 178.2000 133.4000 179.0000 134.6000 ;
	    RECT 182.0000 134.6000 182.8000 139.8000 ;
	    RECT 183.6000 136.0000 184.4000 139.8000 ;
	    RECT 183.6000 135.2000 184.6000 136.0000 ;
	    RECT 182.0000 134.0000 183.2000 134.6000 ;
	    RECT 178.2000 132.6000 182.0000 133.4000 ;
	    RECT 182.6000 132.0000 183.2000 134.0000 ;
	    RECT 182.4000 131.4000 183.2000 132.0000 ;
	    RECT 181.0000 130.8000 181.8000 131.0000 ;
	    RECT 154.8000 130.2000 181.8000 130.8000 ;
	    RECT 154.8000 129.6000 155.6000 130.2000 ;
	    RECT 158.0000 130.0000 159.0000 130.2000 ;
	    RECT 182.4000 129.6000 183.0000 131.4000 ;
	    RECT 183.8000 130.8000 184.6000 135.2000 ;
	    RECT 161.2000 129.4000 162.0000 129.6000 ;
	    RECT 156.6000 129.0000 162.0000 129.4000 ;
	    RECT 155.8000 128.8000 162.0000 129.0000 ;
	    RECT 163.0000 129.0000 171.6000 129.6000 ;
	    RECT 153.2000 128.0000 154.8000 128.8000 ;
	    RECT 155.8000 128.2000 157.2000 128.8000 ;
	    RECT 163.0000 128.2000 163.6000 129.0000 ;
	    RECT 170.8000 128.8000 171.6000 129.0000 ;
	    RECT 174.0000 129.0000 183.0000 129.6000 ;
	    RECT 174.0000 128.8000 174.8000 129.0000 ;
	    RECT 154.2000 127.6000 154.8000 128.0000 ;
	    RECT 157.8000 127.6000 163.6000 128.2000 ;
	    RECT 164.2000 127.6000 166.8000 128.4000 ;
	    RECT 151.6000 126.8000 153.6000 127.4000 ;
	    RECT 154.2000 126.8000 158.4000 127.6000 ;
	    RECT 153.0000 126.2000 153.6000 126.8000 ;
	    RECT 153.0000 125.6000 154.0000 126.2000 ;
	    RECT 153.2000 122.2000 154.0000 125.6000 ;
	    RECT 156.4000 122.2000 157.2000 126.8000 ;
	    RECT 159.6000 122.2000 160.4000 125.0000 ;
	    RECT 161.2000 122.2000 162.0000 125.0000 ;
	    RECT 162.8000 122.2000 163.6000 127.0000 ;
	    RECT 166.0000 122.2000 166.8000 127.0000 ;
	    RECT 169.2000 122.2000 170.0000 128.4000 ;
	    RECT 177.2000 127.6000 179.8000 128.4000 ;
	    RECT 172.4000 126.8000 176.6000 127.6000 ;
	    RECT 170.8000 122.2000 171.6000 125.0000 ;
	    RECT 172.4000 122.2000 173.2000 125.0000 ;
	    RECT 174.0000 122.2000 174.8000 125.0000 ;
	    RECT 177.2000 122.2000 178.0000 127.6000 ;
	    RECT 182.4000 127.4000 183.0000 129.0000 ;
	    RECT 180.4000 126.8000 183.0000 127.4000 ;
	    RECT 183.6000 130.0000 184.6000 130.8000 ;
	    RECT 186.8000 133.8000 187.6000 139.8000 ;
	    RECT 193.2000 136.6000 194.0000 139.8000 ;
	    RECT 194.8000 137.0000 195.6000 139.8000 ;
	    RECT 196.4000 137.0000 197.2000 139.8000 ;
	    RECT 198.0000 137.0000 198.8000 139.8000 ;
	    RECT 201.2000 137.0000 202.0000 139.8000 ;
	    RECT 204.4000 137.0000 205.2000 139.8000 ;
	    RECT 206.0000 137.0000 206.8000 139.8000 ;
	    RECT 207.6000 137.0000 208.4000 139.8000 ;
	    RECT 209.2000 137.0000 210.0000 139.8000 ;
	    RECT 191.4000 135.8000 194.0000 136.6000 ;
	    RECT 210.8000 136.6000 211.6000 139.8000 ;
	    RECT 197.4000 135.8000 202.0000 136.4000 ;
	    RECT 191.4000 135.2000 192.2000 135.8000 ;
	    RECT 189.2000 134.4000 192.2000 135.2000 ;
	    RECT 186.8000 133.0000 195.6000 133.8000 ;
	    RECT 197.4000 133.4000 198.2000 135.8000 ;
	    RECT 201.2000 135.6000 202.0000 135.8000 ;
	    RECT 202.8000 135.6000 204.4000 136.4000 ;
	    RECT 207.4000 135.6000 208.4000 136.4000 ;
	    RECT 210.8000 135.8000 213.2000 136.6000 ;
	    RECT 199.6000 133.6000 200.4000 135.2000 ;
	    RECT 201.2000 134.8000 202.0000 135.0000 ;
	    RECT 201.2000 134.2000 205.6000 134.8000 ;
	    RECT 204.8000 134.0000 205.6000 134.2000 ;
	    RECT 183.6000 128.3000 184.4000 130.0000 ;
	    RECT 185.2000 128.3000 186.0000 128.4000 ;
	    RECT 183.6000 127.7000 186.0000 128.3000 ;
	    RECT 180.4000 122.2000 181.2000 126.8000 ;
	    RECT 183.6000 122.2000 184.4000 127.7000 ;
	    RECT 185.2000 127.6000 186.0000 127.7000 ;
	    RECT 186.8000 127.4000 187.6000 133.0000 ;
	    RECT 196.2000 132.6000 198.2000 133.4000 ;
	    RECT 202.0000 132.6000 205.2000 133.4000 ;
	    RECT 207.6000 132.8000 208.4000 135.6000 ;
	    RECT 212.4000 135.2000 213.2000 135.8000 ;
	    RECT 212.4000 134.6000 214.2000 135.2000 ;
	    RECT 213.4000 133.4000 214.2000 134.6000 ;
	    RECT 217.2000 134.6000 218.0000 139.8000 ;
	    RECT 218.8000 136.0000 219.6000 139.8000 ;
	    RECT 218.8000 135.2000 219.8000 136.0000 ;
	    RECT 217.2000 134.0000 218.4000 134.6000 ;
	    RECT 213.4000 132.6000 217.2000 133.4000 ;
	    RECT 188.2000 132.0000 189.0000 132.2000 ;
	    RECT 190.0000 132.0000 190.8000 132.4000 ;
	    RECT 193.2000 132.0000 194.0000 132.4000 ;
	    RECT 210.8000 132.0000 211.6000 132.6000 ;
	    RECT 217.8000 132.0000 218.4000 134.0000 ;
	    RECT 188.2000 131.4000 211.6000 132.0000 ;
	    RECT 217.6000 131.4000 218.4000 132.0000 ;
	    RECT 217.6000 129.6000 218.2000 131.4000 ;
	    RECT 219.0000 130.8000 219.8000 135.2000 ;
	    RECT 196.4000 129.4000 197.2000 129.6000 ;
	    RECT 191.8000 129.0000 197.2000 129.4000 ;
	    RECT 191.0000 128.8000 197.2000 129.0000 ;
	    RECT 198.2000 129.0000 206.8000 129.6000 ;
	    RECT 188.4000 128.0000 190.0000 128.8000 ;
	    RECT 191.0000 128.2000 192.4000 128.8000 ;
	    RECT 198.2000 128.2000 198.8000 129.0000 ;
	    RECT 206.0000 128.8000 206.8000 129.0000 ;
	    RECT 209.2000 129.0000 218.2000 129.6000 ;
	    RECT 209.2000 128.8000 210.0000 129.0000 ;
	    RECT 189.4000 127.6000 190.0000 128.0000 ;
	    RECT 193.0000 127.6000 198.8000 128.2000 ;
	    RECT 199.4000 127.6000 202.0000 128.4000 ;
	    RECT 186.8000 126.8000 188.8000 127.4000 ;
	    RECT 189.4000 126.8000 193.6000 127.6000 ;
	    RECT 188.2000 126.2000 188.8000 126.8000 ;
	    RECT 188.2000 125.6000 189.2000 126.2000 ;
	    RECT 188.4000 122.2000 189.2000 125.6000 ;
	    RECT 191.6000 122.2000 192.4000 126.8000 ;
	    RECT 194.8000 122.2000 195.6000 125.0000 ;
	    RECT 196.4000 122.2000 197.2000 125.0000 ;
	    RECT 198.0000 122.2000 198.8000 127.0000 ;
	    RECT 201.2000 122.2000 202.0000 127.0000 ;
	    RECT 204.4000 122.2000 205.2000 128.4000 ;
	    RECT 212.4000 127.6000 215.0000 128.4000 ;
	    RECT 207.6000 126.8000 211.8000 127.6000 ;
	    RECT 206.0000 122.2000 206.8000 125.0000 ;
	    RECT 207.6000 122.2000 208.4000 125.0000 ;
	    RECT 209.2000 122.2000 210.0000 125.0000 ;
	    RECT 212.4000 122.2000 213.2000 127.6000 ;
	    RECT 217.6000 127.4000 218.2000 129.0000 ;
	    RECT 215.6000 126.8000 218.2000 127.4000 ;
	    RECT 218.8000 130.0000 219.8000 130.8000 ;
	    RECT 215.6000 122.2000 216.4000 126.8000 ;
	    RECT 218.8000 122.2000 219.6000 130.0000 ;
	    RECT 4.4000 112.4000 5.2000 119.8000 ;
	    RECT 9.2000 112.4000 10.0000 119.8000 ;
	    RECT 3.0000 111.8000 5.2000 112.4000 ;
	    RECT 7.8000 111.8000 10.0000 112.4000 ;
	    RECT 3.0000 111.2000 3.6000 111.8000 ;
	    RECT 7.8000 111.2000 8.4000 111.8000 ;
	    RECT 2.4000 110.4000 3.6000 111.2000 ;
	    RECT 7.2000 110.4000 8.4000 111.2000 ;
	    RECT 3.0000 107.4000 3.6000 110.4000 ;
	    RECT 4.4000 108.8000 5.2000 110.4000 ;
	    RECT 7.8000 107.4000 8.4000 110.4000 ;
	    RECT 9.2000 110.3000 10.0000 110.4000 ;
	    RECT 10.8000 110.3000 11.6000 110.4000 ;
	    RECT 9.2000 109.7000 11.6000 110.3000 ;
	    RECT 9.2000 108.8000 10.0000 109.7000 ;
	    RECT 10.8000 109.6000 11.6000 109.7000 ;
	    RECT 3.0000 106.8000 5.2000 107.4000 ;
	    RECT 7.8000 106.8000 10.0000 107.4000 ;
	    RECT 4.4000 102.2000 5.2000 106.8000 ;
	    RECT 9.2000 102.2000 10.0000 106.8000 ;
	    RECT 10.8000 104.8000 11.6000 106.4000 ;
	    RECT 12.4000 102.2000 13.2000 119.8000 ;
	    RECT 14.0000 114.3000 14.8000 114.4000 ;
	    RECT 15.6000 114.3000 16.4000 119.8000 ;
	    RECT 14.0000 113.7000 16.4000 114.3000 ;
	    RECT 14.0000 113.6000 14.8000 113.7000 ;
	    RECT 15.6000 108.3000 16.4000 113.7000 ;
	    RECT 17.2000 112.4000 18.0000 119.8000 ;
	    RECT 20.4000 112.4000 21.2000 119.8000 ;
	    RECT 17.2000 111.8000 21.2000 112.4000 ;
	    RECT 22.0000 111.8000 22.8000 119.8000 ;
	    RECT 26.2000 112.4000 27.0000 119.8000 ;
	    RECT 27.6000 113.6000 28.4000 114.4000 ;
	    RECT 27.8000 112.4000 28.4000 113.6000 ;
	    RECT 30.0000 112.4000 30.8000 119.8000 ;
	    RECT 33.2000 112.4000 34.0000 119.8000 ;
	    RECT 26.2000 111.8000 27.2000 112.4000 ;
	    RECT 27.8000 111.8000 29.2000 112.4000 ;
	    RECT 30.0000 111.8000 34.0000 112.4000 ;
	    RECT 34.8000 111.8000 35.6000 119.8000 ;
	    RECT 38.0000 112.0000 38.8000 119.8000 ;
	    RECT 41.2000 115.2000 42.0000 119.8000 ;
	    RECT 18.0000 110.4000 18.8000 110.8000 ;
	    RECT 22.0000 110.4000 22.6000 111.8000 ;
	    RECT 17.2000 109.8000 18.8000 110.4000 ;
	    RECT 20.4000 109.8000 22.8000 110.4000 ;
	    RECT 17.2000 109.6000 18.0000 109.8000 ;
	    RECT 18.8000 108.3000 19.6000 109.2000 ;
	    RECT 15.6000 107.7000 19.6000 108.3000 ;
	    RECT 14.0000 104.8000 14.8000 106.4000 ;
	    RECT 15.6000 102.2000 16.4000 107.7000 ;
	    RECT 18.8000 107.6000 19.6000 107.7000 ;
	    RECT 20.4000 106.2000 21.0000 109.8000 ;
	    RECT 22.0000 109.6000 22.8000 109.8000 ;
	    RECT 25.2000 108.8000 26.0000 110.4000 ;
	    RECT 26.6000 108.4000 27.2000 111.8000 ;
	    RECT 28.4000 111.6000 29.2000 111.8000 ;
	    RECT 30.8000 110.4000 31.6000 110.8000 ;
	    RECT 34.8000 110.4000 35.4000 111.8000 ;
	    RECT 37.8000 111.2000 38.8000 112.0000 ;
	    RECT 39.4000 114.6000 42.0000 115.2000 ;
	    RECT 39.4000 113.0000 40.0000 114.6000 ;
	    RECT 44.4000 114.4000 45.2000 119.8000 ;
	    RECT 47.6000 117.0000 48.4000 119.8000 ;
	    RECT 49.2000 117.0000 50.0000 119.8000 ;
	    RECT 50.8000 117.0000 51.6000 119.8000 ;
	    RECT 45.8000 114.4000 50.0000 115.2000 ;
	    RECT 42.6000 113.6000 45.2000 114.4000 ;
	    RECT 52.4000 113.6000 53.2000 119.8000 ;
	    RECT 55.6000 115.0000 56.4000 119.8000 ;
	    RECT 58.8000 115.0000 59.6000 119.8000 ;
	    RECT 60.4000 117.0000 61.2000 119.8000 ;
	    RECT 62.0000 117.0000 62.8000 119.8000 ;
	    RECT 65.2000 115.2000 66.0000 119.8000 ;
	    RECT 68.4000 116.4000 69.2000 119.8000 ;
	    RECT 68.4000 115.8000 69.4000 116.4000 ;
	    RECT 68.8000 115.2000 69.4000 115.8000 ;
	    RECT 64.0000 114.4000 68.2000 115.2000 ;
	    RECT 68.8000 114.6000 70.8000 115.2000 ;
	    RECT 55.6000 113.6000 58.2000 114.4000 ;
	    RECT 58.8000 113.8000 64.6000 114.4000 ;
	    RECT 67.6000 114.0000 68.2000 114.4000 ;
	    RECT 47.6000 113.0000 48.4000 113.2000 ;
	    RECT 39.4000 112.4000 48.4000 113.0000 ;
	    RECT 50.8000 113.0000 51.6000 113.2000 ;
	    RECT 58.8000 113.0000 59.4000 113.8000 ;
	    RECT 65.2000 113.2000 66.6000 113.8000 ;
	    RECT 67.6000 113.2000 69.2000 114.0000 ;
	    RECT 50.8000 112.4000 59.4000 113.0000 ;
	    RECT 60.4000 113.0000 66.6000 113.2000 ;
	    RECT 60.4000 112.6000 65.8000 113.0000 ;
	    RECT 60.4000 112.4000 61.2000 112.6000 ;
	    RECT 30.0000 109.8000 31.6000 110.4000 ;
	    RECT 33.2000 110.3000 35.6000 110.4000 ;
	    RECT 36.4000 110.3000 37.2000 110.4000 ;
	    RECT 33.2000 109.8000 37.2000 110.3000 ;
	    RECT 30.0000 109.6000 30.8000 109.8000 ;
	    RECT 22.0000 108.3000 22.8000 108.4000 ;
	    RECT 23.6000 108.3000 24.4000 108.4000 ;
	    RECT 22.0000 108.2000 24.4000 108.3000 ;
	    RECT 22.0000 107.7000 25.2000 108.2000 ;
	    RECT 22.0000 107.6000 22.8000 107.7000 ;
	    RECT 23.6000 107.6000 25.2000 107.7000 ;
	    RECT 26.6000 107.6000 29.2000 108.4000 ;
	    RECT 31.6000 107.6000 32.4000 109.2000 ;
	    RECT 24.4000 107.2000 25.2000 107.6000 ;
	    RECT 20.4000 102.2000 21.2000 106.2000 ;
	    RECT 22.0000 105.6000 22.8000 106.4000 ;
	    RECT 23.8000 106.2000 27.4000 106.6000 ;
	    RECT 28.4000 106.2000 29.0000 107.6000 ;
	    RECT 33.2000 106.2000 33.8000 109.8000 ;
	    RECT 34.8000 109.7000 37.2000 109.8000 ;
	    RECT 34.8000 109.6000 35.6000 109.7000 ;
	    RECT 36.4000 109.6000 37.2000 109.7000 ;
	    RECT 37.8000 106.8000 38.6000 111.2000 ;
	    RECT 39.4000 110.6000 40.0000 112.4000 ;
	    RECT 39.2000 110.0000 40.0000 110.6000 ;
	    RECT 46.0000 110.0000 69.4000 110.6000 ;
	    RECT 39.2000 108.0000 39.8000 110.0000 ;
	    RECT 46.0000 109.4000 46.8000 110.0000 ;
	    RECT 63.6000 109.6000 64.4000 110.0000 ;
	    RECT 66.8000 109.6000 67.6000 110.0000 ;
	    RECT 68.6000 109.8000 69.4000 110.0000 ;
	    RECT 40.4000 108.6000 44.2000 109.4000 ;
	    RECT 39.2000 107.4000 40.4000 108.0000 ;
	    RECT 23.6000 106.0000 27.6000 106.2000 ;
	    RECT 21.8000 104.8000 22.6000 105.6000 ;
	    RECT 23.6000 102.2000 24.4000 106.0000 ;
	    RECT 26.8000 102.2000 27.6000 106.0000 ;
	    RECT 28.4000 102.2000 29.2000 106.2000 ;
	    RECT 33.2000 102.2000 34.0000 106.2000 ;
	    RECT 34.8000 105.6000 35.6000 106.4000 ;
	    RECT 37.8000 106.0000 38.8000 106.8000 ;
	    RECT 34.6000 104.8000 35.4000 105.6000 ;
	    RECT 38.0000 102.2000 38.8000 106.0000 ;
	    RECT 39.6000 102.2000 40.4000 107.4000 ;
	    RECT 43.4000 107.4000 44.2000 108.6000 ;
	    RECT 43.4000 106.8000 45.2000 107.4000 ;
	    RECT 44.4000 106.2000 45.2000 106.8000 ;
	    RECT 49.2000 106.4000 50.0000 109.2000 ;
	    RECT 52.4000 108.6000 55.6000 109.4000 ;
	    RECT 59.4000 108.6000 61.4000 109.4000 ;
	    RECT 70.0000 109.0000 70.8000 114.6000 ;
	    RECT 52.0000 107.8000 52.8000 108.0000 ;
	    RECT 52.0000 107.2000 56.4000 107.8000 ;
	    RECT 55.6000 107.0000 56.4000 107.2000 ;
	    RECT 57.2000 106.8000 58.0000 108.4000 ;
	    RECT 44.4000 105.4000 46.8000 106.2000 ;
	    RECT 49.2000 105.6000 50.2000 106.4000 ;
	    RECT 53.2000 105.6000 54.8000 106.4000 ;
	    RECT 55.6000 106.2000 56.4000 106.4000 ;
	    RECT 59.4000 106.2000 60.2000 108.6000 ;
	    RECT 62.0000 108.2000 70.8000 109.0000 ;
	    RECT 65.4000 106.8000 68.4000 107.6000 ;
	    RECT 65.4000 106.2000 66.2000 106.8000 ;
	    RECT 55.6000 105.6000 60.2000 106.2000 ;
	    RECT 46.0000 102.2000 46.8000 105.4000 ;
	    RECT 63.6000 105.4000 66.2000 106.2000 ;
	    RECT 47.6000 102.2000 48.4000 105.0000 ;
	    RECT 49.2000 102.2000 50.0000 105.0000 ;
	    RECT 50.8000 102.2000 51.6000 105.0000 ;
	    RECT 52.4000 102.2000 53.2000 105.0000 ;
	    RECT 55.6000 102.2000 56.4000 105.0000 ;
	    RECT 58.8000 102.2000 59.6000 105.0000 ;
	    RECT 60.4000 102.2000 61.2000 105.0000 ;
	    RECT 62.0000 102.2000 62.8000 105.0000 ;
	    RECT 63.6000 102.2000 64.4000 105.4000 ;
	    RECT 70.0000 102.2000 70.8000 108.2000 ;
	    RECT 71.6000 106.3000 72.4000 106.4000 ;
	    RECT 76.4000 106.3000 77.2000 106.4000 ;
	    RECT 71.6000 105.7000 77.2000 106.3000 ;
	    RECT 71.6000 105.6000 72.4000 105.7000 ;
	    RECT 76.4000 104.8000 77.2000 105.7000 ;
	    RECT 78.0000 102.2000 78.8000 119.8000 ;
	    RECT 81.2000 111.2000 82.0000 119.8000 ;
	    RECT 84.4000 111.2000 85.2000 119.8000 ;
	    RECT 87.6000 111.2000 88.4000 119.8000 ;
	    RECT 90.8000 111.2000 91.6000 119.8000 ;
	    RECT 95.6000 116.4000 96.4000 119.8000 ;
	    RECT 95.4000 115.8000 96.4000 116.4000 ;
	    RECT 95.4000 115.2000 96.0000 115.8000 ;
	    RECT 98.8000 115.2000 99.6000 119.8000 ;
	    RECT 102.0000 117.0000 102.8000 119.8000 ;
	    RECT 103.6000 117.0000 104.4000 119.8000 ;
	    RECT 79.6000 110.4000 82.0000 111.2000 ;
	    RECT 83.0000 110.4000 85.2000 111.2000 ;
	    RECT 86.2000 110.4000 88.4000 111.2000 ;
	    RECT 89.8000 110.4000 91.6000 111.2000 ;
	    RECT 94.0000 114.6000 96.0000 115.2000 ;
	    RECT 79.6000 107.6000 80.4000 110.4000 ;
	    RECT 83.0000 109.0000 83.8000 110.4000 ;
	    RECT 86.2000 109.0000 87.0000 110.4000 ;
	    RECT 89.8000 109.0000 90.6000 110.4000 ;
	    RECT 81.2000 108.2000 83.8000 109.0000 ;
	    RECT 84.6000 108.2000 87.0000 109.0000 ;
	    RECT 88.0000 108.2000 90.6000 109.0000 ;
	    RECT 83.0000 107.6000 83.8000 108.2000 ;
	    RECT 86.2000 107.6000 87.0000 108.2000 ;
	    RECT 89.8000 107.6000 90.6000 108.2000 ;
	    RECT 94.0000 109.0000 94.8000 114.6000 ;
	    RECT 96.6000 114.4000 100.8000 115.2000 ;
	    RECT 105.2000 115.0000 106.0000 119.8000 ;
	    RECT 108.4000 115.0000 109.2000 119.8000 ;
	    RECT 96.6000 114.0000 97.2000 114.4000 ;
	    RECT 95.6000 113.2000 97.2000 114.0000 ;
	    RECT 100.2000 113.8000 106.0000 114.4000 ;
	    RECT 98.2000 113.2000 99.6000 113.8000 ;
	    RECT 98.2000 113.0000 104.4000 113.2000 ;
	    RECT 99.0000 112.6000 104.4000 113.0000 ;
	    RECT 103.6000 112.4000 104.4000 112.6000 ;
	    RECT 105.4000 113.0000 106.0000 113.8000 ;
	    RECT 106.6000 113.6000 109.2000 114.4000 ;
	    RECT 111.6000 113.6000 112.4000 119.8000 ;
	    RECT 113.2000 117.0000 114.0000 119.8000 ;
	    RECT 114.8000 117.0000 115.6000 119.8000 ;
	    RECT 116.4000 117.0000 117.2000 119.8000 ;
	    RECT 114.8000 114.4000 119.0000 115.2000 ;
	    RECT 119.6000 114.4000 120.4000 119.8000 ;
	    RECT 122.8000 115.2000 123.6000 119.8000 ;
	    RECT 122.8000 114.6000 125.4000 115.2000 ;
	    RECT 119.6000 113.6000 122.2000 114.4000 ;
	    RECT 113.2000 113.0000 114.0000 113.2000 ;
	    RECT 105.4000 112.4000 114.0000 113.0000 ;
	    RECT 116.4000 113.0000 117.2000 113.2000 ;
	    RECT 124.8000 113.0000 125.4000 114.6000 ;
	    RECT 116.4000 112.4000 125.4000 113.0000 ;
	    RECT 124.8000 110.6000 125.4000 112.4000 ;
	    RECT 126.0000 112.0000 126.8000 119.8000 ;
	    RECT 130.8000 115.8000 131.6000 119.8000 ;
	    RECT 131.0000 115.6000 131.6000 115.8000 ;
	    RECT 134.0000 115.8000 134.8000 119.8000 ;
	    RECT 134.0000 115.6000 134.6000 115.8000 ;
	    RECT 131.0000 115.0000 134.6000 115.6000 ;
	    RECT 132.4000 112.8000 133.2000 114.4000 ;
	    RECT 134.0000 112.4000 134.6000 115.0000 ;
	    RECT 126.0000 111.2000 127.0000 112.0000 ;
	    RECT 95.4000 110.0000 118.8000 110.6000 ;
	    RECT 124.8000 110.0000 125.6000 110.6000 ;
	    RECT 95.4000 109.8000 96.2000 110.0000 ;
	    RECT 98.8000 109.6000 99.6000 110.0000 ;
	    RECT 100.4000 109.6000 101.2000 110.0000 ;
	    RECT 118.0000 109.4000 118.8000 110.0000 ;
	    RECT 94.0000 108.2000 102.8000 109.0000 ;
	    RECT 103.4000 108.6000 105.4000 109.4000 ;
	    RECT 109.2000 108.6000 112.4000 109.4000 ;
	    RECT 79.6000 106.8000 82.0000 107.6000 ;
	    RECT 83.0000 106.8000 85.2000 107.6000 ;
	    RECT 86.2000 106.8000 88.4000 107.6000 ;
	    RECT 89.8000 106.8000 91.6000 107.6000 ;
	    RECT 81.2000 102.2000 82.0000 106.8000 ;
	    RECT 84.4000 102.2000 85.2000 106.8000 ;
	    RECT 87.6000 102.2000 88.4000 106.8000 ;
	    RECT 90.8000 102.2000 91.6000 106.8000 ;
	    RECT 94.0000 102.2000 94.8000 108.2000 ;
	    RECT 96.4000 106.8000 99.4000 107.6000 ;
	    RECT 98.6000 106.2000 99.4000 106.8000 ;
	    RECT 104.6000 106.2000 105.4000 108.6000 ;
	    RECT 106.8000 106.8000 107.6000 108.4000 ;
	    RECT 112.0000 107.8000 112.8000 108.0000 ;
	    RECT 108.4000 107.2000 112.8000 107.8000 ;
	    RECT 108.4000 107.0000 109.2000 107.2000 ;
	    RECT 114.8000 106.4000 115.6000 109.2000 ;
	    RECT 120.6000 108.6000 124.4000 109.4000 ;
	    RECT 120.6000 107.4000 121.4000 108.6000 ;
	    RECT 125.0000 108.0000 125.6000 110.0000 ;
	    RECT 108.4000 106.2000 109.2000 106.4000 ;
	    RECT 98.6000 105.4000 101.2000 106.2000 ;
	    RECT 104.6000 105.6000 109.2000 106.2000 ;
	    RECT 110.0000 105.6000 111.6000 106.4000 ;
	    RECT 114.6000 105.6000 115.6000 106.4000 ;
	    RECT 119.6000 106.8000 121.4000 107.4000 ;
	    RECT 124.4000 107.4000 125.6000 108.0000 ;
	    RECT 126.2000 110.3000 127.0000 111.2000 ;
	    RECT 129.2000 110.3000 130.0000 112.4000 ;
	    RECT 134.0000 111.6000 134.8000 112.4000 ;
	    RECT 126.2000 109.7000 130.0000 110.3000 ;
	    RECT 119.6000 106.2000 120.4000 106.8000 ;
	    RECT 100.4000 102.2000 101.2000 105.4000 ;
	    RECT 118.0000 105.4000 120.4000 106.2000 ;
	    RECT 102.0000 102.2000 102.8000 105.0000 ;
	    RECT 103.6000 102.2000 104.4000 105.0000 ;
	    RECT 105.2000 102.2000 106.0000 105.0000 ;
	    RECT 108.4000 102.2000 109.2000 105.0000 ;
	    RECT 111.6000 102.2000 112.4000 105.0000 ;
	    RECT 113.2000 102.2000 114.0000 105.0000 ;
	    RECT 114.8000 102.2000 115.6000 105.0000 ;
	    RECT 116.4000 102.2000 117.2000 105.0000 ;
	    RECT 118.0000 102.2000 118.8000 105.4000 ;
	    RECT 124.4000 102.2000 125.2000 107.4000 ;
	    RECT 126.2000 106.8000 127.0000 109.7000 ;
	    RECT 130.8000 109.6000 132.4000 110.4000 ;
	    RECT 134.0000 108.4000 134.6000 111.6000 ;
	    RECT 133.0000 108.2000 134.6000 108.4000 ;
	    RECT 126.0000 106.0000 127.0000 106.8000 ;
	    RECT 132.8000 107.8000 134.6000 108.2000 ;
	    RECT 137.2000 110.3000 138.0000 119.8000 ;
	    RECT 141.4000 112.6000 142.2000 119.8000 ;
	    RECT 140.4000 111.8000 142.2000 112.6000 ;
	    RECT 140.4000 111.6000 141.2000 111.8000 ;
	    RECT 138.8000 110.3000 139.6000 110.4000 ;
	    RECT 137.2000 109.7000 139.6000 110.3000 ;
	    RECT 126.0000 102.2000 126.8000 106.0000 ;
	    RECT 132.8000 102.2000 133.6000 107.8000 ;
	    RECT 135.6000 104.8000 136.4000 106.4000 ;
	    RECT 137.2000 102.2000 138.0000 109.7000 ;
	    RECT 138.8000 109.6000 139.6000 109.7000 ;
	    RECT 140.6000 108.4000 141.2000 111.6000 ;
	    RECT 142.0000 109.6000 142.8000 111.2000 ;
	    RECT 140.4000 107.6000 141.2000 108.4000 ;
	    RECT 138.8000 104.8000 139.6000 106.4000 ;
	    RECT 140.6000 104.2000 141.2000 107.6000 ;
	    RECT 140.4000 102.2000 141.2000 104.2000 ;
	    RECT 143.6000 102.2000 144.4000 119.8000 ;
	    RECT 149.0000 114.4000 149.8000 119.8000 ;
	    RECT 147.6000 113.6000 148.4000 114.4000 ;
	    RECT 149.0000 113.6000 150.8000 114.4000 ;
	    RECT 147.6000 112.4000 148.2000 113.6000 ;
	    RECT 149.0000 112.4000 149.8000 113.6000 ;
	    RECT 155.8000 112.6000 156.6000 119.8000 ;
	    RECT 146.8000 111.8000 148.2000 112.4000 ;
	    RECT 148.8000 111.8000 149.8000 112.4000 ;
	    RECT 154.8000 111.8000 156.6000 112.6000 ;
	    RECT 162.8000 112.4000 163.6000 119.8000 ;
	    RECT 166.0000 112.4000 166.8000 119.8000 ;
	    RECT 162.8000 111.8000 166.8000 112.4000 ;
	    RECT 167.6000 111.8000 168.4000 119.8000 ;
	    RECT 171.8000 112.4000 172.6000 119.8000 ;
	    RECT 175.6000 119.2000 179.6000 119.8000 ;
	    RECT 173.2000 113.6000 174.0000 114.4000 ;
	    RECT 173.4000 112.4000 174.0000 113.6000 ;
	    RECT 171.8000 111.8000 172.8000 112.4000 ;
	    RECT 173.4000 111.8000 174.8000 112.4000 ;
	    RECT 175.6000 111.8000 176.4000 119.2000 ;
	    RECT 177.2000 111.8000 178.0000 118.6000 ;
	    RECT 178.8000 112.4000 179.6000 119.2000 ;
	    RECT 182.0000 112.4000 182.8000 119.8000 ;
	    RECT 178.8000 111.8000 182.8000 112.4000 ;
	    RECT 146.8000 111.6000 147.6000 111.8000 ;
	    RECT 148.8000 108.4000 149.4000 111.8000 ;
	    RECT 150.0000 108.8000 150.8000 110.4000 ;
	    RECT 155.0000 108.4000 155.6000 111.8000 ;
	    RECT 156.4000 109.6000 157.2000 111.2000 ;
	    RECT 163.6000 110.4000 164.4000 110.8000 ;
	    RECT 167.6000 110.4000 168.2000 111.8000 ;
	    RECT 162.8000 110.3000 164.4000 110.4000 ;
	    RECT 159.7000 109.8000 164.4000 110.3000 ;
	    RECT 166.0000 109.8000 168.4000 110.4000 ;
	    RECT 159.7000 109.7000 163.6000 109.8000 ;
	    RECT 146.8000 107.6000 149.4000 108.4000 ;
	    RECT 151.6000 108.3000 152.4000 108.4000 ;
	    RECT 154.8000 108.3000 155.6000 108.4000 ;
	    RECT 159.7000 108.3000 160.3000 109.7000 ;
	    RECT 162.8000 109.6000 163.6000 109.7000 ;
	    RECT 151.6000 108.2000 160.3000 108.3000 ;
	    RECT 150.8000 107.7000 160.3000 108.2000 ;
	    RECT 150.8000 107.6000 152.4000 107.7000 ;
	    RECT 154.8000 107.6000 155.6000 107.7000 ;
	    RECT 164.4000 107.6000 165.2000 109.2000 ;
	    RECT 145.2000 104.8000 146.0000 106.4000 ;
	    RECT 147.0000 106.2000 147.6000 107.6000 ;
	    RECT 150.8000 107.2000 151.6000 107.6000 ;
	    RECT 148.6000 106.2000 152.2000 106.6000 ;
	    RECT 146.8000 102.2000 147.6000 106.2000 ;
	    RECT 148.4000 106.0000 152.4000 106.2000 ;
	    RECT 148.4000 102.2000 149.2000 106.0000 ;
	    RECT 151.6000 102.2000 152.4000 106.0000 ;
	    RECT 153.2000 104.8000 154.0000 106.4000 ;
	    RECT 155.0000 104.2000 155.6000 107.6000 ;
	    RECT 154.8000 102.2000 155.6000 104.2000 ;
	    RECT 166.0000 106.2000 166.6000 109.8000 ;
	    RECT 167.6000 109.6000 168.4000 109.8000 ;
	    RECT 170.8000 108.8000 171.6000 110.4000 ;
	    RECT 172.2000 110.3000 172.8000 111.8000 ;
	    RECT 174.0000 111.6000 174.8000 111.8000 ;
	    RECT 177.4000 111.2000 178.0000 111.8000 ;
	    RECT 175.6000 110.3000 176.4000 111.2000 ;
	    RECT 177.4000 110.6000 179.4000 111.2000 ;
	    RECT 172.2000 109.7000 176.4000 110.3000 ;
	    RECT 172.2000 108.4000 172.8000 109.7000 ;
	    RECT 175.6000 109.6000 176.4000 109.7000 ;
	    RECT 178.8000 110.4000 179.4000 110.6000 ;
	    RECT 181.2000 110.4000 182.0000 110.8000 ;
	    RECT 178.8000 109.6000 179.6000 110.4000 ;
	    RECT 181.2000 109.8000 182.8000 110.4000 ;
	    RECT 182.0000 109.6000 182.8000 109.8000 ;
	    RECT 177.4000 108.8000 178.2000 109.6000 ;
	    RECT 177.4000 108.4000 178.0000 108.8000 ;
	    RECT 169.2000 108.2000 170.0000 108.4000 ;
	    RECT 169.2000 107.6000 170.8000 108.2000 ;
	    RECT 172.2000 107.6000 174.8000 108.4000 ;
	    RECT 175.6000 108.3000 176.4000 108.4000 ;
	    RECT 177.2000 108.3000 178.0000 108.4000 ;
	    RECT 175.6000 107.7000 178.0000 108.3000 ;
	    RECT 175.6000 107.6000 176.4000 107.7000 ;
	    RECT 177.2000 107.6000 178.0000 107.7000 ;
	    RECT 170.0000 107.2000 170.8000 107.6000 ;
	    RECT 166.0000 102.2000 166.8000 106.2000 ;
	    RECT 167.6000 105.6000 168.4000 106.4000 ;
	    RECT 169.4000 106.2000 173.0000 106.6000 ;
	    RECT 174.0000 106.2000 174.6000 107.6000 ;
	    RECT 178.8000 106.2000 179.4000 109.6000 ;
	    RECT 180.4000 107.6000 181.2000 109.2000 ;
	    RECT 169.2000 106.0000 173.2000 106.2000 ;
	    RECT 167.4000 104.8000 168.2000 105.6000 ;
	    RECT 169.2000 102.2000 170.0000 106.0000 ;
	    RECT 172.4000 102.2000 173.2000 106.0000 ;
	    RECT 174.0000 102.2000 174.8000 106.2000 ;
	    RECT 178.2000 104.4000 179.8000 106.2000 ;
	    RECT 177.2000 103.6000 179.8000 104.4000 ;
	    RECT 178.2000 102.2000 179.8000 103.6000 ;
	    RECT 183.6000 102.2000 184.4000 119.8000 ;
	    RECT 186.8000 112.4000 187.6000 119.8000 ;
	    RECT 193.8000 118.4000 194.6000 119.8000 ;
	    RECT 193.8000 117.6000 195.6000 118.4000 ;
	    RECT 192.4000 113.6000 193.2000 114.4000 ;
	    RECT 192.4000 112.4000 193.0000 113.6000 ;
	    RECT 193.8000 112.4000 194.6000 117.6000 ;
	    RECT 198.8000 113.6000 199.6000 114.4000 ;
	    RECT 198.8000 112.4000 199.4000 113.6000 ;
	    RECT 200.2000 112.4000 201.0000 119.8000 ;
	    RECT 186.8000 111.8000 189.0000 112.4000 ;
	    RECT 188.4000 111.2000 189.0000 111.8000 ;
	    RECT 191.6000 111.8000 193.0000 112.4000 ;
	    RECT 193.6000 111.8000 194.6000 112.4000 ;
	    RECT 198.0000 111.8000 199.4000 112.4000 ;
	    RECT 200.0000 111.8000 201.0000 112.4000 ;
	    RECT 191.6000 111.6000 192.4000 111.8000 ;
	    RECT 188.4000 110.4000 189.6000 111.2000 ;
	    RECT 186.8000 108.8000 187.6000 110.4000 ;
	    RECT 188.4000 107.4000 189.0000 110.4000 ;
	    RECT 193.6000 108.4000 194.2000 111.8000 ;
	    RECT 198.0000 111.6000 198.8000 111.8000 ;
	    RECT 194.8000 110.3000 195.6000 110.4000 ;
	    RECT 200.0000 110.3000 200.6000 111.8000 ;
	    RECT 194.8000 109.7000 200.6000 110.3000 ;
	    RECT 194.8000 108.8000 195.6000 109.7000 ;
	    RECT 200.0000 108.4000 200.6000 109.7000 ;
	    RECT 201.2000 110.3000 202.0000 110.4000 ;
	    RECT 206.0000 110.3000 206.8000 119.8000 ;
	    RECT 207.6000 111.6000 208.4000 113.2000 ;
	    RECT 209.2000 112.4000 210.0000 119.8000 ;
	    RECT 212.4000 112.4000 213.2000 119.8000 ;
	    RECT 209.2000 111.8000 213.2000 112.4000 ;
	    RECT 214.0000 111.8000 214.8000 119.8000 ;
	    RECT 201.2000 109.7000 206.8000 110.3000 ;
	    RECT 207.7000 110.3000 208.3000 111.6000 ;
	    RECT 210.0000 110.4000 210.8000 110.8000 ;
	    RECT 214.0000 110.4000 214.6000 111.8000 ;
	    RECT 209.2000 110.3000 210.8000 110.4000 ;
	    RECT 207.7000 109.8000 210.8000 110.3000 ;
	    RECT 212.4000 109.8000 214.8000 110.4000 ;
	    RECT 207.7000 109.7000 210.0000 109.8000 ;
	    RECT 201.2000 108.8000 202.0000 109.7000 ;
	    RECT 191.6000 107.6000 194.2000 108.4000 ;
	    RECT 196.4000 108.2000 197.2000 108.4000 ;
	    RECT 195.6000 107.6000 197.2000 108.2000 ;
	    RECT 198.0000 107.6000 200.6000 108.4000 ;
	    RECT 186.8000 106.8000 189.0000 107.4000 ;
	    RECT 185.2000 104.8000 186.0000 106.4000 ;
	    RECT 186.8000 102.2000 187.6000 106.8000 ;
	    RECT 191.8000 106.2000 192.4000 107.6000 ;
	    RECT 195.6000 107.2000 196.4000 107.6000 ;
	    RECT 193.4000 106.2000 197.0000 106.6000 ;
	    RECT 198.2000 106.2000 198.8000 107.6000 ;
	    RECT 204.4000 106.8000 205.2000 108.4000 ;
	    RECT 199.8000 106.2000 203.4000 106.6000 ;
	    RECT 206.0000 106.2000 206.8000 109.7000 ;
	    RECT 209.2000 109.6000 210.0000 109.7000 ;
	    RECT 210.8000 107.6000 211.6000 109.2000 ;
	    RECT 212.4000 106.2000 213.0000 109.8000 ;
	    RECT 214.0000 109.6000 214.8000 109.8000 ;
	    RECT 214.0000 106.3000 214.8000 106.4000 ;
	    RECT 215.6000 106.3000 216.4000 119.8000 ;
	    RECT 218.8000 112.4000 219.6000 119.8000 ;
	    RECT 218.8000 111.8000 221.0000 112.4000 ;
	    RECT 220.4000 111.2000 221.0000 111.8000 ;
	    RECT 220.4000 110.4000 221.6000 111.2000 ;
	    RECT 218.8000 108.8000 219.6000 110.4000 ;
	    RECT 220.4000 107.4000 221.0000 110.4000 ;
	    RECT 191.6000 102.2000 192.4000 106.2000 ;
	    RECT 193.2000 106.0000 197.2000 106.2000 ;
	    RECT 193.2000 102.2000 194.0000 106.0000 ;
	    RECT 196.4000 102.2000 197.2000 106.0000 ;
	    RECT 198.0000 102.2000 198.8000 106.2000 ;
	    RECT 199.6000 106.0000 203.6000 106.2000 ;
	    RECT 199.6000 102.2000 200.4000 106.0000 ;
	    RECT 202.8000 102.2000 203.6000 106.0000 ;
	    RECT 206.0000 105.6000 207.8000 106.2000 ;
	    RECT 207.0000 104.4000 207.8000 105.6000 ;
	    RECT 207.0000 103.6000 208.4000 104.4000 ;
	    RECT 207.0000 102.2000 207.8000 103.6000 ;
	    RECT 212.4000 102.2000 213.2000 106.2000 ;
	    RECT 214.0000 105.7000 216.4000 106.3000 ;
	    RECT 214.0000 105.6000 214.8000 105.7000 ;
	    RECT 213.8000 104.8000 214.6000 105.6000 ;
	    RECT 215.6000 102.2000 216.4000 105.7000 ;
	    RECT 218.8000 106.8000 221.0000 107.4000 ;
	    RECT 218.8000 102.2000 219.6000 106.8000 ;
	    RECT 2.8000 96.0000 3.6000 99.8000 ;
	    RECT 2.6000 95.2000 3.6000 96.0000 ;
	    RECT 2.6000 90.8000 3.4000 95.2000 ;
	    RECT 4.4000 94.6000 5.2000 99.8000 ;
	    RECT 10.8000 96.6000 11.6000 99.8000 ;
	    RECT 12.4000 97.0000 13.2000 99.8000 ;
	    RECT 14.0000 97.0000 14.8000 99.8000 ;
	    RECT 15.6000 97.0000 16.4000 99.8000 ;
	    RECT 17.2000 97.0000 18.0000 99.8000 ;
	    RECT 20.4000 97.0000 21.2000 99.8000 ;
	    RECT 23.6000 97.0000 24.4000 99.8000 ;
	    RECT 25.2000 97.0000 26.0000 99.8000 ;
	    RECT 26.8000 97.0000 27.6000 99.8000 ;
	    RECT 9.2000 95.8000 11.6000 96.6000 ;
	    RECT 28.4000 96.6000 29.2000 99.8000 ;
	    RECT 9.2000 95.2000 10.0000 95.8000 ;
	    RECT 4.0000 94.0000 5.2000 94.6000 ;
	    RECT 8.2000 94.6000 10.0000 95.2000 ;
	    RECT 14.0000 95.6000 15.0000 96.4000 ;
	    RECT 18.0000 95.6000 19.6000 96.4000 ;
	    RECT 20.4000 95.8000 25.0000 96.4000 ;
	    RECT 28.4000 95.8000 31.0000 96.6000 ;
	    RECT 20.4000 95.6000 21.2000 95.8000 ;
	    RECT 4.0000 92.0000 4.6000 94.0000 ;
	    RECT 8.2000 93.4000 9.0000 94.6000 ;
	    RECT 5.2000 92.6000 9.0000 93.4000 ;
	    RECT 14.0000 92.8000 14.8000 95.6000 ;
	    RECT 20.4000 94.8000 21.2000 95.0000 ;
	    RECT 16.8000 94.2000 21.2000 94.8000 ;
	    RECT 16.8000 94.0000 17.6000 94.2000 ;
	    RECT 22.0000 93.6000 22.8000 95.2000 ;
	    RECT 24.2000 93.4000 25.0000 95.8000 ;
	    RECT 30.2000 95.2000 31.0000 95.8000 ;
	    RECT 30.2000 94.4000 33.2000 95.2000 ;
	    RECT 34.8000 93.8000 35.6000 99.8000 ;
	    RECT 39.6000 95.2000 40.4000 99.8000 ;
	    RECT 41.2000 95.8000 42.0000 99.8000 ;
	    RECT 42.8000 96.0000 43.6000 99.8000 ;
	    RECT 46.0000 96.0000 46.8000 99.8000 ;
	    RECT 42.8000 95.8000 46.8000 96.0000 ;
	    RECT 47.6000 95.8000 48.4000 99.8000 ;
	    RECT 52.0000 96.2000 53.6000 99.8000 ;
	    RECT 17.2000 92.6000 20.4000 93.4000 ;
	    RECT 24.2000 92.6000 26.2000 93.4000 ;
	    RECT 26.8000 93.0000 35.6000 93.8000 ;
	    RECT 10.8000 92.0000 11.6000 92.6000 ;
	    RECT 28.4000 92.0000 29.2000 92.4000 ;
	    RECT 30.0000 92.0000 30.8000 92.4000 ;
	    RECT 33.4000 92.0000 34.2000 92.2000 ;
	    RECT 4.0000 91.4000 4.8000 92.0000 ;
	    RECT 10.8000 91.4000 34.2000 92.0000 ;
	    RECT 2.6000 90.0000 3.6000 90.8000 ;
	    RECT 2.8000 82.2000 3.6000 90.0000 ;
	    RECT 4.2000 89.6000 4.8000 91.4000 ;
	    RECT 4.2000 89.0000 13.2000 89.6000 ;
	    RECT 4.2000 87.4000 4.8000 89.0000 ;
	    RECT 12.4000 88.8000 13.2000 89.0000 ;
	    RECT 15.6000 89.0000 24.2000 89.6000 ;
	    RECT 15.6000 88.8000 16.4000 89.0000 ;
	    RECT 7.4000 87.6000 10.0000 88.4000 ;
	    RECT 4.2000 86.8000 6.8000 87.4000 ;
	    RECT 6.0000 82.2000 6.8000 86.8000 ;
	    RECT 9.2000 82.2000 10.0000 87.6000 ;
	    RECT 10.6000 86.8000 14.8000 87.6000 ;
	    RECT 12.4000 82.2000 13.2000 85.0000 ;
	    RECT 14.0000 82.2000 14.8000 85.0000 ;
	    RECT 15.6000 82.2000 16.4000 85.0000 ;
	    RECT 17.2000 82.2000 18.0000 88.4000 ;
	    RECT 20.4000 87.6000 23.0000 88.4000 ;
	    RECT 23.6000 88.2000 24.2000 89.0000 ;
	    RECT 25.2000 89.4000 26.0000 89.6000 ;
	    RECT 25.2000 89.0000 30.6000 89.4000 ;
	    RECT 25.2000 88.8000 31.4000 89.0000 ;
	    RECT 30.0000 88.2000 31.4000 88.8000 ;
	    RECT 23.6000 87.6000 29.4000 88.2000 ;
	    RECT 32.4000 88.0000 34.0000 88.8000 ;
	    RECT 32.4000 87.6000 33.0000 88.0000 ;
	    RECT 20.4000 82.2000 21.2000 87.0000 ;
	    RECT 23.6000 82.2000 24.4000 87.0000 ;
	    RECT 28.8000 86.8000 33.0000 87.6000 ;
	    RECT 34.8000 87.4000 35.6000 93.0000 ;
	    RECT 38.2000 94.6000 40.4000 95.2000 ;
	    RECT 38.2000 91.6000 38.8000 94.6000 ;
	    RECT 41.4000 94.4000 42.0000 95.8000 ;
	    RECT 43.0000 95.4000 46.6000 95.8000 ;
	    RECT 47.6000 95.2000 50.0000 95.8000 ;
	    RECT 49.2000 95.0000 50.0000 95.2000 ;
	    RECT 50.6000 94.8000 51.4000 95.6000 ;
	    RECT 45.2000 94.4000 46.0000 94.8000 ;
	    RECT 50.6000 94.4000 51.2000 94.8000 ;
	    RECT 41.2000 93.6000 43.8000 94.4000 ;
	    RECT 45.2000 93.8000 46.8000 94.4000 ;
	    RECT 46.0000 93.6000 46.8000 93.8000 ;
	    RECT 47.6000 93.6000 49.2000 94.4000 ;
	    RECT 50.4000 93.6000 51.2000 94.4000 ;
	    RECT 39.6000 91.6000 40.4000 93.2000 ;
	    RECT 37.6000 90.8000 38.8000 91.6000 ;
	    RECT 38.2000 90.2000 38.8000 90.8000 ;
	    RECT 41.2000 90.2000 42.0000 90.4000 ;
	    RECT 43.2000 90.2000 43.8000 93.6000 ;
	    RECT 44.4000 91.6000 45.2000 93.2000 ;
	    RECT 52.0000 92.8000 52.6000 96.2000 ;
	    RECT 57.2000 95.8000 58.0000 99.8000 ;
	    RECT 53.2000 95.4000 54.8000 95.6000 ;
	    RECT 53.2000 94.8000 55.2000 95.4000 ;
	    RECT 55.8000 95.2000 58.0000 95.8000 ;
	    RECT 55.8000 95.0000 56.6000 95.2000 ;
	    RECT 54.6000 94.4000 55.2000 94.8000 ;
	    RECT 53.2000 93.4000 54.0000 94.2000 ;
	    RECT 54.6000 93.8000 58.0000 94.4000 ;
	    RECT 56.4000 93.6000 58.0000 93.8000 ;
	    RECT 51.6000 92.4000 52.6000 92.8000 ;
	    RECT 50.8000 92.2000 52.6000 92.4000 ;
	    RECT 53.4000 92.8000 54.0000 93.4000 ;
	    RECT 53.4000 92.2000 56.0000 92.8000 ;
	    RECT 50.8000 91.6000 52.2000 92.2000 ;
	    RECT 55.2000 92.0000 56.0000 92.2000 ;
	    RECT 58.8000 92.4000 59.6000 99.8000 ;
	    RECT 62.0000 95.2000 62.8000 99.8000 ;
	    RECT 70.0000 96.0000 70.8000 99.8000 ;
	    RECT 60.6000 94.6000 62.8000 95.2000 ;
	    RECT 69.8000 95.2000 70.8000 96.0000 ;
	    RECT 51.6000 90.2000 52.2000 91.6000 ;
	    RECT 53.0000 91.4000 53.8000 91.6000 ;
	    RECT 53.0000 90.8000 56.4000 91.4000 ;
	    RECT 55.8000 90.2000 56.4000 90.8000 ;
	    RECT 58.8000 90.2000 59.4000 92.4000 ;
	    RECT 60.6000 91.6000 61.2000 94.6000 ;
	    RECT 62.0000 92.3000 62.8000 93.2000 ;
	    RECT 68.4000 92.3000 69.2000 92.4000 ;
	    RECT 62.0000 91.7000 69.2000 92.3000 ;
	    RECT 62.0000 91.6000 62.8000 91.7000 ;
	    RECT 68.4000 91.6000 69.2000 91.7000 ;
	    RECT 60.0000 90.8000 61.2000 91.6000 ;
	    RECT 60.6000 90.2000 61.2000 90.8000 ;
	    RECT 69.8000 90.8000 70.6000 95.2000 ;
	    RECT 71.6000 94.6000 72.4000 99.8000 ;
	    RECT 78.0000 96.6000 78.8000 99.8000 ;
	    RECT 79.6000 97.0000 80.4000 99.8000 ;
	    RECT 81.2000 97.0000 82.0000 99.8000 ;
	    RECT 82.8000 97.0000 83.6000 99.8000 ;
	    RECT 84.4000 97.0000 85.2000 99.8000 ;
	    RECT 87.6000 97.0000 88.4000 99.8000 ;
	    RECT 90.8000 97.0000 91.6000 99.8000 ;
	    RECT 92.4000 97.0000 93.2000 99.8000 ;
	    RECT 94.0000 97.0000 94.8000 99.8000 ;
	    RECT 76.4000 95.8000 78.8000 96.6000 ;
	    RECT 95.6000 96.6000 96.4000 99.8000 ;
	    RECT 76.4000 95.2000 77.2000 95.8000 ;
	    RECT 71.2000 94.0000 72.4000 94.6000 ;
	    RECT 75.4000 94.6000 77.2000 95.2000 ;
	    RECT 81.2000 95.6000 82.2000 96.4000 ;
	    RECT 85.2000 95.6000 86.8000 96.4000 ;
	    RECT 87.6000 95.8000 92.2000 96.4000 ;
	    RECT 95.6000 95.8000 98.2000 96.6000 ;
	    RECT 87.6000 95.6000 88.4000 95.8000 ;
	    RECT 71.2000 92.0000 71.8000 94.0000 ;
	    RECT 75.4000 93.4000 76.2000 94.6000 ;
	    RECT 72.4000 92.6000 76.2000 93.4000 ;
	    RECT 81.2000 92.8000 82.0000 95.6000 ;
	    RECT 87.6000 94.8000 88.4000 95.0000 ;
	    RECT 84.0000 94.2000 88.4000 94.8000 ;
	    RECT 84.0000 94.0000 84.8000 94.2000 ;
	    RECT 89.2000 93.6000 90.0000 95.2000 ;
	    RECT 91.4000 93.4000 92.2000 95.8000 ;
	    RECT 97.4000 95.2000 98.2000 95.8000 ;
	    RECT 97.4000 94.4000 100.4000 95.2000 ;
	    RECT 102.0000 93.8000 102.8000 99.8000 ;
	    RECT 84.4000 92.6000 87.6000 93.4000 ;
	    RECT 91.4000 92.6000 93.4000 93.4000 ;
	    RECT 94.0000 93.0000 102.8000 93.8000 ;
	    RECT 78.0000 92.0000 78.8000 92.6000 ;
	    RECT 95.6000 92.0000 96.4000 92.4000 ;
	    RECT 98.8000 92.0000 99.6000 92.4000 ;
	    RECT 100.6000 92.0000 101.4000 92.2000 ;
	    RECT 71.2000 91.4000 72.0000 92.0000 ;
	    RECT 78.0000 91.4000 101.4000 92.0000 ;
	    RECT 38.2000 89.6000 40.4000 90.2000 ;
	    RECT 41.2000 89.6000 42.6000 90.2000 ;
	    RECT 43.2000 89.6000 44.2000 90.2000 ;
	    RECT 33.6000 86.8000 35.6000 87.4000 ;
	    RECT 25.2000 82.2000 26.0000 85.0000 ;
	    RECT 26.8000 82.2000 27.6000 85.0000 ;
	    RECT 30.0000 82.2000 30.8000 86.8000 ;
	    RECT 33.6000 86.2000 34.2000 86.8000 ;
	    RECT 33.2000 85.6000 34.2000 86.2000 ;
	    RECT 33.2000 82.2000 34.0000 85.6000 ;
	    RECT 39.6000 82.2000 40.4000 89.6000 ;
	    RECT 42.0000 88.4000 42.6000 89.6000 ;
	    RECT 42.0000 87.6000 42.8000 88.4000 ;
	    RECT 43.4000 82.2000 44.2000 89.6000 ;
	    RECT 47.6000 89.6000 50.0000 90.2000 ;
	    RECT 51.6000 89.6000 53.6000 90.2000 ;
	    RECT 47.6000 82.2000 48.4000 89.6000 ;
	    RECT 49.2000 89.4000 50.0000 89.6000 ;
	    RECT 52.0000 84.4000 53.6000 89.6000 ;
	    RECT 55.8000 89.6000 58.0000 90.2000 ;
	    RECT 55.8000 89.4000 56.6000 89.6000 ;
	    RECT 50.8000 83.6000 53.6000 84.4000 ;
	    RECT 52.0000 82.2000 53.6000 83.6000 ;
	    RECT 57.2000 82.2000 58.0000 89.6000 ;
	    RECT 58.8000 82.2000 59.6000 90.2000 ;
	    RECT 60.6000 89.6000 62.8000 90.2000 ;
	    RECT 69.8000 90.0000 70.8000 90.8000 ;
	    RECT 62.0000 82.2000 62.8000 89.6000 ;
	    RECT 70.0000 82.2000 70.8000 90.0000 ;
	    RECT 71.4000 89.6000 72.0000 91.4000 ;
	    RECT 71.4000 89.0000 80.4000 89.6000 ;
	    RECT 71.4000 87.4000 72.0000 89.0000 ;
	    RECT 79.6000 88.8000 80.4000 89.0000 ;
	    RECT 82.8000 89.0000 91.4000 89.6000 ;
	    RECT 82.8000 88.8000 83.6000 89.0000 ;
	    RECT 74.6000 87.6000 77.2000 88.4000 ;
	    RECT 71.4000 86.8000 74.0000 87.4000 ;
	    RECT 73.2000 82.2000 74.0000 86.8000 ;
	    RECT 76.4000 82.2000 77.2000 87.6000 ;
	    RECT 77.8000 86.8000 82.0000 87.6000 ;
	    RECT 79.6000 82.2000 80.4000 85.0000 ;
	    RECT 81.2000 82.2000 82.0000 85.0000 ;
	    RECT 82.8000 82.2000 83.6000 85.0000 ;
	    RECT 84.4000 82.2000 85.2000 88.4000 ;
	    RECT 87.6000 87.6000 90.2000 88.4000 ;
	    RECT 90.8000 88.2000 91.4000 89.0000 ;
	    RECT 92.4000 89.4000 93.2000 89.6000 ;
	    RECT 92.4000 89.0000 97.8000 89.4000 ;
	    RECT 92.4000 88.8000 98.6000 89.0000 ;
	    RECT 97.2000 88.2000 98.6000 88.8000 ;
	    RECT 90.8000 87.6000 96.6000 88.2000 ;
	    RECT 99.6000 88.0000 101.2000 88.8000 ;
	    RECT 99.6000 87.6000 100.2000 88.0000 ;
	    RECT 87.6000 82.2000 88.4000 87.0000 ;
	    RECT 90.8000 82.2000 91.6000 87.0000 ;
	    RECT 96.0000 86.8000 100.2000 87.6000 ;
	    RECT 102.0000 87.4000 102.8000 93.0000 ;
	    RECT 100.8000 86.8000 102.8000 87.4000 ;
	    RECT 103.6000 92.4000 104.4000 99.8000 ;
	    RECT 106.8000 95.2000 107.6000 99.8000 ;
	    RECT 105.4000 94.6000 107.6000 95.2000 ;
	    RECT 103.6000 90.2000 104.2000 92.4000 ;
	    RECT 105.4000 91.6000 106.0000 94.6000 ;
	    RECT 106.8000 91.6000 107.6000 93.2000 ;
	    RECT 108.4000 92.4000 109.2000 99.8000 ;
	    RECT 111.6000 95.2000 112.4000 99.8000 ;
	    RECT 110.2000 94.6000 112.4000 95.2000 ;
	    RECT 113.2000 95.2000 114.0000 99.8000 ;
	    RECT 113.2000 94.6000 115.4000 95.2000 ;
	    RECT 104.8000 90.8000 106.0000 91.6000 ;
	    RECT 105.4000 90.2000 106.0000 90.8000 ;
	    RECT 108.4000 90.2000 109.0000 92.4000 ;
	    RECT 110.2000 91.6000 110.8000 94.6000 ;
	    RECT 111.6000 92.3000 112.4000 93.2000 ;
	    RECT 113.2000 92.3000 114.0000 93.2000 ;
	    RECT 111.6000 91.7000 114.0000 92.3000 ;
	    RECT 111.6000 91.6000 112.4000 91.7000 ;
	    RECT 113.2000 91.6000 114.0000 91.7000 ;
	    RECT 114.8000 91.6000 115.4000 94.6000 ;
	    RECT 116.4000 92.4000 117.2000 99.8000 ;
	    RECT 119.2000 94.2000 120.0000 99.8000 ;
	    RECT 109.6000 90.8000 110.8000 91.6000 ;
	    RECT 110.2000 90.2000 110.8000 90.8000 ;
	    RECT 114.8000 90.8000 116.0000 91.6000 ;
	    RECT 114.8000 90.2000 115.4000 90.8000 ;
	    RECT 116.6000 90.2000 117.2000 92.4000 ;
	    RECT 118.2000 93.8000 120.0000 94.2000 ;
	    RECT 128.0000 94.2000 128.8000 99.8000 ;
	    RECT 128.0000 93.8000 129.8000 94.2000 ;
	    RECT 118.2000 93.6000 119.8000 93.8000 ;
	    RECT 128.2000 93.6000 129.8000 93.8000 ;
	    RECT 118.2000 90.4000 118.8000 93.6000 ;
	    RECT 120.4000 91.6000 122.0000 92.4000 ;
	    RECT 126.0000 91.6000 127.6000 92.4000 ;
	    RECT 92.4000 82.2000 93.2000 85.0000 ;
	    RECT 94.0000 82.2000 94.8000 85.0000 ;
	    RECT 97.2000 82.2000 98.0000 86.8000 ;
	    RECT 100.8000 86.2000 101.4000 86.8000 ;
	    RECT 100.4000 85.6000 101.4000 86.2000 ;
	    RECT 100.4000 82.2000 101.2000 85.6000 ;
	    RECT 103.6000 82.2000 104.4000 90.2000 ;
	    RECT 105.4000 89.6000 107.6000 90.2000 ;
	    RECT 106.8000 82.2000 107.6000 89.6000 ;
	    RECT 108.4000 82.2000 109.2000 90.2000 ;
	    RECT 110.2000 89.6000 112.4000 90.2000 ;
	    RECT 111.6000 82.2000 112.4000 89.6000 ;
	    RECT 113.2000 89.6000 115.4000 90.2000 ;
	    RECT 113.2000 82.2000 114.0000 89.6000 ;
	    RECT 116.4000 82.2000 117.2000 90.2000 ;
	    RECT 118.0000 89.6000 118.8000 90.4000 ;
	    RECT 122.8000 90.3000 123.6000 91.2000 ;
	    RECT 124.4000 90.3000 125.2000 91.2000 ;
	    RECT 122.8000 89.7000 125.2000 90.3000 ;
	    RECT 122.8000 89.6000 123.6000 89.7000 ;
	    RECT 124.4000 89.6000 125.2000 89.7000 ;
	    RECT 129.2000 90.4000 129.8000 93.6000 ;
	    RECT 129.2000 89.6000 130.0000 90.4000 ;
	    RECT 118.2000 87.0000 118.8000 89.6000 ;
	    RECT 119.6000 87.6000 120.4000 89.2000 ;
	    RECT 127.6000 87.6000 128.4000 89.2000 ;
	    RECT 129.2000 87.0000 129.8000 89.6000 ;
	    RECT 118.2000 86.4000 121.8000 87.0000 ;
	    RECT 118.2000 86.2000 118.8000 86.4000 ;
	    RECT 118.0000 82.2000 118.8000 86.2000 ;
	    RECT 121.2000 86.2000 121.8000 86.4000 ;
	    RECT 126.2000 86.4000 129.8000 87.0000 ;
	    RECT 126.2000 86.2000 126.8000 86.4000 ;
	    RECT 121.2000 82.2000 122.0000 86.2000 ;
	    RECT 126.0000 82.2000 126.8000 86.2000 ;
	    RECT 129.2000 86.2000 129.8000 86.4000 ;
	    RECT 129.2000 82.2000 130.0000 86.2000 ;
	    RECT 130.8000 82.2000 131.6000 99.8000 ;
	    RECT 132.4000 95.6000 133.2000 97.2000 ;
	    RECT 135.6000 96.0000 136.4000 99.8000 ;
	    RECT 135.4000 95.2000 136.4000 96.0000 ;
	    RECT 135.4000 90.8000 136.2000 95.2000 ;
	    RECT 137.2000 94.6000 138.0000 99.8000 ;
	    RECT 143.6000 96.6000 144.4000 99.8000 ;
	    RECT 145.2000 97.0000 146.0000 99.8000 ;
	    RECT 146.8000 97.0000 147.6000 99.8000 ;
	    RECT 148.4000 97.0000 149.2000 99.8000 ;
	    RECT 150.0000 97.0000 150.8000 99.8000 ;
	    RECT 153.2000 97.0000 154.0000 99.8000 ;
	    RECT 156.4000 97.0000 157.2000 99.8000 ;
	    RECT 158.0000 97.0000 158.8000 99.8000 ;
	    RECT 159.6000 97.0000 160.4000 99.8000 ;
	    RECT 142.0000 95.8000 144.4000 96.6000 ;
	    RECT 161.2000 96.6000 162.0000 99.8000 ;
	    RECT 142.0000 95.2000 142.8000 95.8000 ;
	    RECT 136.8000 94.0000 138.0000 94.6000 ;
	    RECT 141.0000 94.6000 142.8000 95.2000 ;
	    RECT 146.8000 95.6000 147.8000 96.4000 ;
	    RECT 150.8000 95.6000 152.4000 96.4000 ;
	    RECT 153.2000 95.8000 157.8000 96.4000 ;
	    RECT 161.2000 95.8000 163.8000 96.6000 ;
	    RECT 153.2000 95.6000 154.0000 95.8000 ;
	    RECT 136.8000 92.0000 137.4000 94.0000 ;
	    RECT 141.0000 93.4000 141.8000 94.6000 ;
	    RECT 138.0000 92.6000 141.8000 93.4000 ;
	    RECT 146.8000 92.8000 147.6000 95.6000 ;
	    RECT 153.2000 94.8000 154.0000 95.0000 ;
	    RECT 149.6000 94.2000 154.0000 94.8000 ;
	    RECT 149.6000 94.0000 150.4000 94.2000 ;
	    RECT 154.8000 93.6000 155.6000 95.2000 ;
	    RECT 157.0000 93.4000 157.8000 95.8000 ;
	    RECT 163.0000 95.2000 163.8000 95.8000 ;
	    RECT 163.0000 94.4000 166.0000 95.2000 ;
	    RECT 167.6000 93.8000 168.4000 99.8000 ;
	    RECT 150.0000 92.6000 153.2000 93.4000 ;
	    RECT 157.0000 92.6000 159.0000 93.4000 ;
	    RECT 159.6000 93.0000 168.4000 93.8000 ;
	    RECT 143.6000 92.0000 144.4000 92.6000 ;
	    RECT 161.2000 92.0000 162.0000 92.4000 ;
	    RECT 166.2000 92.0000 167.0000 92.2000 ;
	    RECT 136.8000 91.4000 137.6000 92.0000 ;
	    RECT 143.6000 91.4000 167.0000 92.0000 ;
	    RECT 135.4000 90.0000 136.4000 90.8000 ;
	    RECT 135.6000 82.2000 136.4000 90.0000 ;
	    RECT 137.0000 89.6000 137.6000 91.4000 ;
	    RECT 137.0000 89.0000 146.0000 89.6000 ;
	    RECT 137.0000 87.4000 137.6000 89.0000 ;
	    RECT 145.2000 88.8000 146.0000 89.0000 ;
	    RECT 148.4000 89.0000 157.0000 89.6000 ;
	    RECT 148.4000 88.8000 149.2000 89.0000 ;
	    RECT 140.2000 87.6000 142.8000 88.4000 ;
	    RECT 137.0000 86.8000 139.6000 87.4000 ;
	    RECT 138.8000 82.2000 139.6000 86.8000 ;
	    RECT 142.0000 82.2000 142.8000 87.6000 ;
	    RECT 143.4000 86.8000 147.6000 87.6000 ;
	    RECT 145.2000 82.2000 146.0000 85.0000 ;
	    RECT 146.8000 82.2000 147.6000 85.0000 ;
	    RECT 148.4000 82.2000 149.2000 85.0000 ;
	    RECT 150.0000 82.2000 150.8000 88.4000 ;
	    RECT 153.2000 87.6000 155.8000 88.4000 ;
	    RECT 156.4000 88.2000 157.0000 89.0000 ;
	    RECT 158.0000 89.4000 158.8000 89.6000 ;
	    RECT 158.0000 89.0000 163.4000 89.4000 ;
	    RECT 158.0000 88.8000 164.2000 89.0000 ;
	    RECT 162.8000 88.2000 164.2000 88.8000 ;
	    RECT 156.4000 87.6000 162.2000 88.2000 ;
	    RECT 165.2000 88.0000 166.8000 88.8000 ;
	    RECT 165.2000 87.6000 165.8000 88.0000 ;
	    RECT 153.2000 82.2000 154.0000 87.0000 ;
	    RECT 156.4000 82.2000 157.2000 87.0000 ;
	    RECT 161.6000 86.8000 165.8000 87.6000 ;
	    RECT 167.6000 87.4000 168.4000 93.0000 ;
	    RECT 166.4000 86.8000 168.4000 87.4000 ;
	    RECT 174.0000 93.8000 174.8000 99.8000 ;
	    RECT 180.4000 96.6000 181.2000 99.8000 ;
	    RECT 182.0000 97.0000 182.8000 99.8000 ;
	    RECT 183.6000 97.0000 184.4000 99.8000 ;
	    RECT 185.2000 97.0000 186.0000 99.8000 ;
	    RECT 188.4000 97.0000 189.2000 99.8000 ;
	    RECT 191.6000 97.0000 192.4000 99.8000 ;
	    RECT 193.2000 97.0000 194.0000 99.8000 ;
	    RECT 194.8000 97.0000 195.6000 99.8000 ;
	    RECT 196.4000 97.0000 197.2000 99.8000 ;
	    RECT 178.6000 95.8000 181.2000 96.6000 ;
	    RECT 198.0000 96.6000 198.8000 99.8000 ;
	    RECT 184.6000 95.8000 189.2000 96.4000 ;
	    RECT 178.6000 95.2000 179.4000 95.8000 ;
	    RECT 176.4000 94.4000 179.4000 95.2000 ;
	    RECT 174.0000 93.0000 182.8000 93.8000 ;
	    RECT 184.6000 93.4000 185.4000 95.8000 ;
	    RECT 188.4000 95.6000 189.2000 95.8000 ;
	    RECT 190.0000 95.6000 191.6000 96.4000 ;
	    RECT 194.6000 95.6000 195.6000 96.4000 ;
	    RECT 198.0000 95.8000 200.4000 96.6000 ;
	    RECT 186.8000 93.6000 187.6000 95.2000 ;
	    RECT 188.4000 94.8000 189.2000 95.0000 ;
	    RECT 188.4000 94.2000 192.8000 94.8000 ;
	    RECT 192.0000 94.0000 192.8000 94.2000 ;
	    RECT 174.0000 87.4000 174.8000 93.0000 ;
	    RECT 183.4000 92.6000 185.4000 93.4000 ;
	    RECT 189.2000 92.6000 192.4000 93.4000 ;
	    RECT 194.8000 92.8000 195.6000 95.6000 ;
	    RECT 199.6000 95.2000 200.4000 95.8000 ;
	    RECT 199.6000 94.6000 201.4000 95.2000 ;
	    RECT 200.6000 93.4000 201.4000 94.6000 ;
	    RECT 204.4000 94.6000 205.2000 99.8000 ;
	    RECT 206.0000 96.0000 206.8000 99.8000 ;
	    RECT 209.8000 98.4000 210.6000 99.8000 ;
	    RECT 209.2000 97.6000 210.6000 98.4000 ;
	    RECT 209.8000 96.4000 210.6000 97.6000 ;
	    RECT 206.0000 95.2000 207.0000 96.0000 ;
	    RECT 209.8000 95.8000 211.6000 96.4000 ;
	    RECT 214.0000 96.0000 214.8000 99.8000 ;
	    RECT 217.2000 96.0000 218.0000 99.8000 ;
	    RECT 214.0000 95.8000 218.0000 96.0000 ;
	    RECT 218.8000 95.8000 219.6000 99.8000 ;
	    RECT 204.4000 94.0000 205.6000 94.6000 ;
	    RECT 200.6000 92.6000 204.4000 93.4000 ;
	    RECT 175.4000 92.0000 176.2000 92.2000 ;
	    RECT 177.2000 92.0000 178.0000 92.4000 ;
	    RECT 180.4000 92.0000 181.2000 92.4000 ;
	    RECT 198.0000 92.0000 198.8000 92.6000 ;
	    RECT 205.0000 92.0000 205.6000 94.0000 ;
	    RECT 175.4000 91.4000 198.8000 92.0000 ;
	    RECT 204.8000 91.4000 205.6000 92.0000 ;
	    RECT 204.8000 89.6000 205.4000 91.4000 ;
	    RECT 206.2000 90.8000 207.0000 95.2000 ;
	    RECT 183.6000 89.4000 184.4000 89.6000 ;
	    RECT 179.0000 89.0000 184.4000 89.4000 ;
	    RECT 178.2000 88.8000 184.4000 89.0000 ;
	    RECT 185.4000 89.0000 194.0000 89.6000 ;
	    RECT 175.6000 88.0000 177.2000 88.8000 ;
	    RECT 178.2000 88.2000 179.6000 88.8000 ;
	    RECT 185.4000 88.2000 186.0000 89.0000 ;
	    RECT 193.2000 88.8000 194.0000 89.0000 ;
	    RECT 196.4000 89.0000 205.4000 89.6000 ;
	    RECT 196.4000 88.8000 197.2000 89.0000 ;
	    RECT 176.6000 87.6000 177.2000 88.0000 ;
	    RECT 180.2000 87.6000 186.0000 88.2000 ;
	    RECT 186.6000 87.6000 189.2000 88.4000 ;
	    RECT 174.0000 86.8000 176.0000 87.4000 ;
	    RECT 176.6000 86.8000 180.8000 87.6000 ;
	    RECT 158.0000 82.2000 158.8000 85.0000 ;
	    RECT 159.6000 82.2000 160.4000 85.0000 ;
	    RECT 162.8000 82.2000 163.6000 86.8000 ;
	    RECT 166.4000 86.2000 167.0000 86.8000 ;
	    RECT 166.0000 85.6000 167.0000 86.2000 ;
	    RECT 175.4000 86.2000 176.0000 86.8000 ;
	    RECT 175.4000 85.6000 176.4000 86.2000 ;
	    RECT 166.0000 82.2000 166.8000 85.6000 ;
	    RECT 175.6000 82.2000 176.4000 85.6000 ;
	    RECT 178.8000 82.2000 179.6000 86.8000 ;
	    RECT 182.0000 82.2000 182.8000 85.0000 ;
	    RECT 183.6000 82.2000 184.4000 85.0000 ;
	    RECT 185.2000 82.2000 186.0000 87.0000 ;
	    RECT 188.4000 82.2000 189.2000 87.0000 ;
	    RECT 191.6000 82.2000 192.4000 88.4000 ;
	    RECT 199.6000 87.6000 202.2000 88.4000 ;
	    RECT 194.8000 86.8000 199.0000 87.6000 ;
	    RECT 193.2000 82.2000 194.0000 85.0000 ;
	    RECT 194.8000 82.2000 195.6000 85.0000 ;
	    RECT 196.4000 82.2000 197.2000 85.0000 ;
	    RECT 199.6000 82.2000 200.4000 87.6000 ;
	    RECT 204.8000 87.4000 205.4000 89.0000 ;
	    RECT 202.8000 86.8000 205.4000 87.4000 ;
	    RECT 206.0000 90.0000 207.0000 90.8000 ;
	    RECT 202.8000 82.2000 203.6000 86.8000 ;
	    RECT 206.0000 82.2000 206.8000 90.0000 ;
	    RECT 209.2000 88.8000 210.0000 90.4000 ;
	    RECT 210.8000 82.2000 211.6000 95.8000 ;
	    RECT 214.2000 95.4000 217.8000 95.8000 ;
	    RECT 212.4000 93.6000 213.2000 95.2000 ;
	    RECT 218.8000 94.4000 219.4000 95.8000 ;
	    RECT 217.0000 93.6000 219.6000 94.4000 ;
	    RECT 224.0000 94.2000 224.8000 99.8000 ;
	    RECT 224.0000 93.8000 225.8000 94.2000 ;
	    RECT 224.2000 93.6000 225.8000 93.8000 ;
	    RECT 215.6000 91.6000 216.4000 93.2000 ;
	    RECT 217.0000 90.4000 217.6000 93.6000 ;
	    RECT 222.0000 91.6000 223.6000 92.4000 ;
	    RECT 215.6000 89.6000 217.6000 90.4000 ;
	    RECT 220.4000 89.6000 221.2000 91.2000 ;
	    RECT 225.2000 90.4000 225.8000 93.6000 ;
	    RECT 225.2000 89.6000 226.0000 90.4000 ;
	    RECT 216.6000 82.2000 217.4000 89.6000 ;
	    RECT 223.6000 87.6000 224.4000 89.2000 ;
	    RECT 225.2000 87.0000 225.8000 89.6000 ;
	    RECT 222.2000 86.4000 225.8000 87.0000 ;
	    RECT 222.0000 82.2000 222.8000 86.4000 ;
	    RECT 225.2000 86.2000 225.8000 86.4000 ;
	    RECT 225.2000 82.2000 226.0000 86.2000 ;
	    RECT 2.8000 72.0000 3.6000 79.8000 ;
	    RECT 6.0000 75.2000 6.8000 79.8000 ;
	    RECT 2.6000 71.2000 3.6000 72.0000 ;
	    RECT 4.2000 74.6000 6.8000 75.2000 ;
	    RECT 4.2000 73.0000 4.8000 74.6000 ;
	    RECT 9.2000 74.4000 10.0000 79.8000 ;
	    RECT 12.4000 77.0000 13.2000 79.8000 ;
	    RECT 14.0000 77.0000 14.8000 79.8000 ;
	    RECT 15.6000 77.0000 16.4000 79.8000 ;
	    RECT 10.6000 74.4000 14.8000 75.2000 ;
	    RECT 7.4000 73.6000 10.0000 74.4000 ;
	    RECT 17.2000 73.6000 18.0000 79.8000 ;
	    RECT 20.4000 75.0000 21.2000 79.8000 ;
	    RECT 23.6000 75.0000 24.4000 79.8000 ;
	    RECT 25.2000 77.0000 26.0000 79.8000 ;
	    RECT 26.8000 77.0000 27.6000 79.8000 ;
	    RECT 30.0000 75.2000 30.8000 79.8000 ;
	    RECT 33.2000 76.4000 34.0000 79.8000 ;
	    RECT 33.2000 75.8000 34.2000 76.4000 ;
	    RECT 33.6000 75.2000 34.2000 75.8000 ;
	    RECT 28.8000 74.4000 33.0000 75.2000 ;
	    RECT 33.6000 74.6000 35.6000 75.2000 ;
	    RECT 20.4000 73.6000 23.0000 74.4000 ;
	    RECT 23.6000 73.8000 29.4000 74.4000 ;
	    RECT 32.4000 74.0000 33.0000 74.4000 ;
	    RECT 12.4000 73.0000 13.2000 73.2000 ;
	    RECT 4.2000 72.4000 13.2000 73.0000 ;
	    RECT 15.6000 73.0000 16.4000 73.2000 ;
	    RECT 23.6000 73.0000 24.2000 73.8000 ;
	    RECT 30.0000 73.2000 31.4000 73.8000 ;
	    RECT 32.4000 73.2000 34.0000 74.0000 ;
	    RECT 15.6000 72.4000 24.2000 73.0000 ;
	    RECT 25.2000 73.0000 31.4000 73.2000 ;
	    RECT 25.2000 72.6000 30.6000 73.0000 ;
	    RECT 25.2000 72.4000 26.0000 72.6000 ;
	    RECT 2.6000 66.8000 3.4000 71.2000 ;
	    RECT 4.2000 70.6000 4.8000 72.4000 ;
	    RECT 4.0000 70.0000 4.8000 70.6000 ;
	    RECT 10.8000 70.0000 34.2000 70.6000 ;
	    RECT 4.0000 68.0000 4.6000 70.0000 ;
	    RECT 10.8000 69.4000 11.6000 70.0000 ;
	    RECT 28.4000 69.6000 29.2000 70.0000 ;
	    RECT 30.0000 69.6000 30.8000 70.0000 ;
	    RECT 31.6000 69.6000 32.4000 70.0000 ;
	    RECT 33.4000 69.8000 34.2000 70.0000 ;
	    RECT 5.2000 68.6000 9.0000 69.4000 ;
	    RECT 4.0000 67.4000 5.2000 68.0000 ;
	    RECT 2.6000 66.0000 3.6000 66.8000 ;
	    RECT 2.8000 62.2000 3.6000 66.0000 ;
	    RECT 4.4000 62.2000 5.2000 67.4000 ;
	    RECT 8.2000 67.4000 9.0000 68.6000 ;
	    RECT 8.2000 66.8000 10.0000 67.4000 ;
	    RECT 9.2000 66.2000 10.0000 66.8000 ;
	    RECT 14.0000 66.4000 14.8000 69.2000 ;
	    RECT 17.2000 68.6000 20.4000 69.4000 ;
	    RECT 24.2000 68.6000 26.2000 69.4000 ;
	    RECT 34.8000 69.0000 35.6000 74.6000 ;
	    RECT 39.0000 72.4000 39.8000 79.8000 ;
	    RECT 40.4000 73.6000 42.0000 74.4000 ;
	    RECT 43.6000 73.6000 44.4000 74.4000 ;
	    RECT 40.6000 72.4000 41.2000 73.6000 ;
	    RECT 43.6000 72.4000 44.2000 73.6000 ;
	    RECT 45.0000 72.4000 45.8000 79.8000 ;
	    RECT 39.0000 71.8000 40.0000 72.4000 ;
	    RECT 40.6000 72.3000 42.0000 72.4000 ;
	    RECT 42.8000 72.3000 44.2000 72.4000 ;
	    RECT 40.6000 71.8000 44.2000 72.3000 ;
	    RECT 44.8000 71.8000 45.8000 72.4000 ;
	    RECT 49.2000 72.4000 50.0000 79.8000 ;
	    RECT 52.4000 72.4000 53.2000 79.8000 ;
	    RECT 49.2000 71.8000 53.2000 72.4000 ;
	    RECT 16.8000 67.8000 17.6000 68.0000 ;
	    RECT 16.8000 67.2000 21.2000 67.8000 ;
	    RECT 20.4000 67.0000 21.2000 67.2000 ;
	    RECT 22.0000 66.8000 22.8000 68.4000 ;
	    RECT 9.2000 65.4000 11.6000 66.2000 ;
	    RECT 14.0000 65.6000 15.0000 66.4000 ;
	    RECT 18.0000 65.6000 19.6000 66.4000 ;
	    RECT 20.4000 66.2000 21.2000 66.4000 ;
	    RECT 24.2000 66.2000 25.0000 68.6000 ;
	    RECT 26.8000 68.2000 35.6000 69.0000 ;
	    RECT 38.0000 68.8000 38.8000 70.4000 ;
	    RECT 39.4000 68.4000 40.0000 71.8000 ;
	    RECT 41.2000 71.7000 43.6000 71.8000 ;
	    RECT 41.2000 71.6000 42.0000 71.7000 ;
	    RECT 42.8000 71.6000 43.6000 71.7000 ;
	    RECT 44.8000 68.4000 45.4000 71.8000 ;
	    RECT 54.0000 71.6000 54.8000 79.8000 ;
	    RECT 58.2000 72.4000 59.0000 79.8000 ;
	    RECT 59.6000 73.6000 60.4000 74.4000 ;
	    RECT 59.8000 72.4000 60.4000 73.6000 ;
	    RECT 58.2000 71.8000 59.2000 72.4000 ;
	    RECT 59.8000 72.3000 61.2000 72.4000 ;
	    RECT 66.8000 72.3000 67.6000 72.4000 ;
	    RECT 59.8000 71.8000 67.6000 72.3000 ;
	    RECT 50.0000 70.4000 50.8000 70.8000 ;
	    RECT 54.0000 70.4000 54.6000 71.6000 ;
	    RECT 46.0000 68.8000 46.8000 70.4000 ;
	    RECT 49.2000 69.8000 50.8000 70.4000 ;
	    RECT 52.4000 69.8000 54.8000 70.4000 ;
	    RECT 49.2000 69.6000 50.0000 69.8000 ;
	    RECT 30.2000 66.8000 33.2000 67.6000 ;
	    RECT 30.2000 66.2000 31.0000 66.8000 ;
	    RECT 20.4000 65.6000 25.0000 66.2000 ;
	    RECT 10.8000 62.2000 11.6000 65.4000 ;
	    RECT 28.4000 65.4000 31.0000 66.2000 ;
	    RECT 12.4000 62.2000 13.2000 65.0000 ;
	    RECT 14.0000 62.2000 14.8000 65.0000 ;
	    RECT 15.6000 62.2000 16.4000 65.0000 ;
	    RECT 17.2000 62.2000 18.0000 65.0000 ;
	    RECT 20.4000 62.2000 21.2000 65.0000 ;
	    RECT 23.6000 62.2000 24.4000 65.0000 ;
	    RECT 25.2000 62.2000 26.0000 65.0000 ;
	    RECT 26.8000 62.2000 27.6000 65.0000 ;
	    RECT 28.4000 62.2000 29.2000 65.4000 ;
	    RECT 34.8000 62.2000 35.6000 68.2000 ;
	    RECT 36.4000 68.2000 37.2000 68.4000 ;
	    RECT 36.4000 67.6000 38.0000 68.2000 ;
	    RECT 39.4000 67.6000 42.0000 68.4000 ;
	    RECT 42.8000 67.6000 45.4000 68.4000 ;
	    RECT 47.6000 68.2000 48.4000 68.4000 ;
	    RECT 46.8000 67.6000 48.4000 68.2000 ;
	    RECT 50.8000 67.6000 51.6000 69.2000 ;
	    RECT 37.2000 67.2000 38.0000 67.6000 ;
	    RECT 36.6000 66.2000 40.2000 66.6000 ;
	    RECT 41.2000 66.2000 41.8000 67.6000 ;
	    RECT 43.0000 66.2000 43.6000 67.6000 ;
	    RECT 46.8000 67.2000 47.6000 67.6000 ;
	    RECT 44.6000 66.2000 48.2000 66.6000 ;
	    RECT 52.4000 66.2000 53.0000 69.8000 ;
	    RECT 54.0000 69.6000 54.8000 69.8000 ;
	    RECT 57.2000 68.8000 58.0000 70.4000 ;
	    RECT 58.6000 68.4000 59.2000 71.8000 ;
	    RECT 60.4000 71.7000 67.6000 71.8000 ;
	    RECT 60.4000 71.6000 61.2000 71.7000 ;
	    RECT 66.8000 71.6000 67.6000 71.7000 ;
	    RECT 55.6000 68.2000 56.4000 68.4000 ;
	    RECT 55.6000 67.6000 57.2000 68.2000 ;
	    RECT 58.6000 67.6000 61.2000 68.4000 ;
	    RECT 56.4000 67.2000 57.2000 67.6000 ;
	    RECT 36.4000 66.0000 40.4000 66.2000 ;
	    RECT 36.4000 62.2000 37.2000 66.0000 ;
	    RECT 39.6000 62.2000 40.4000 66.0000 ;
	    RECT 41.2000 62.2000 42.0000 66.2000 ;
	    RECT 42.8000 62.2000 43.6000 66.2000 ;
	    RECT 44.4000 66.0000 48.4000 66.2000 ;
	    RECT 44.4000 62.2000 45.2000 66.0000 ;
	    RECT 47.6000 62.2000 48.4000 66.0000 ;
	    RECT 52.4000 62.2000 53.2000 66.2000 ;
	    RECT 54.0000 65.6000 54.8000 66.4000 ;
	    RECT 55.8000 66.2000 59.4000 66.6000 ;
	    RECT 60.4000 66.2000 61.0000 67.6000 ;
	    RECT 55.6000 66.0000 59.6000 66.2000 ;
	    RECT 53.8000 64.8000 54.6000 65.6000 ;
	    RECT 55.6000 62.2000 56.4000 66.0000 ;
	    RECT 58.8000 62.2000 59.6000 66.0000 ;
	    RECT 60.4000 62.2000 61.2000 66.2000 ;
	    RECT 66.8000 64.8000 67.6000 66.4000 ;
	    RECT 68.4000 62.2000 69.2000 79.8000 ;
	    RECT 70.6000 72.6000 71.4000 79.8000 ;
	    RECT 75.6000 73.6000 76.4000 74.4000 ;
	    RECT 70.6000 71.8000 72.4000 72.6000 ;
	    RECT 75.6000 72.4000 76.2000 73.6000 ;
	    RECT 77.0000 72.4000 77.8000 79.8000 ;
	    RECT 82.8000 76.4000 83.6000 79.8000 ;
	    RECT 82.6000 75.8000 83.6000 76.4000 ;
	    RECT 82.6000 75.2000 83.2000 75.8000 ;
	    RECT 86.0000 75.2000 86.8000 79.8000 ;
	    RECT 89.2000 77.0000 90.0000 79.8000 ;
	    RECT 90.8000 77.0000 91.6000 79.8000 ;
	    RECT 74.8000 71.8000 76.2000 72.4000 ;
	    RECT 76.8000 71.8000 77.8000 72.4000 ;
	    RECT 81.2000 74.6000 83.2000 75.2000 ;
	    RECT 70.0000 69.6000 70.8000 71.2000 ;
	    RECT 71.6000 68.4000 72.2000 71.8000 ;
	    RECT 74.8000 71.6000 75.6000 71.8000 ;
	    RECT 76.8000 68.4000 77.4000 71.8000 ;
	    RECT 78.0000 68.8000 78.8000 70.4000 ;
	    RECT 81.2000 69.0000 82.0000 74.6000 ;
	    RECT 83.8000 74.4000 88.0000 75.2000 ;
	    RECT 92.4000 75.0000 93.2000 79.8000 ;
	    RECT 95.6000 75.0000 96.4000 79.8000 ;
	    RECT 83.8000 74.0000 84.4000 74.4000 ;
	    RECT 82.8000 73.2000 84.4000 74.0000 ;
	    RECT 87.4000 73.8000 93.2000 74.4000 ;
	    RECT 85.4000 73.2000 86.8000 73.8000 ;
	    RECT 85.4000 73.0000 91.6000 73.2000 ;
	    RECT 86.2000 72.6000 91.6000 73.0000 ;
	    RECT 90.8000 72.4000 91.6000 72.6000 ;
	    RECT 92.6000 73.0000 93.2000 73.8000 ;
	    RECT 93.8000 73.6000 96.4000 74.4000 ;
	    RECT 98.8000 73.6000 99.6000 79.8000 ;
	    RECT 100.4000 77.0000 101.2000 79.8000 ;
	    RECT 102.0000 77.0000 102.8000 79.8000 ;
	    RECT 103.6000 77.0000 104.4000 79.8000 ;
	    RECT 102.0000 74.4000 106.2000 75.2000 ;
	    RECT 106.8000 74.4000 107.6000 79.8000 ;
	    RECT 110.0000 75.2000 110.8000 79.8000 ;
	    RECT 110.0000 74.6000 112.6000 75.2000 ;
	    RECT 106.8000 73.6000 109.4000 74.4000 ;
	    RECT 100.4000 73.0000 101.2000 73.2000 ;
	    RECT 92.6000 72.4000 101.2000 73.0000 ;
	    RECT 103.6000 73.0000 104.4000 73.2000 ;
	    RECT 112.0000 73.0000 112.6000 74.6000 ;
	    RECT 103.6000 72.4000 112.6000 73.0000 ;
	    RECT 112.0000 70.6000 112.6000 72.4000 ;
	    RECT 113.2000 72.0000 114.0000 79.8000 ;
	    RECT 113.2000 71.2000 114.2000 72.0000 ;
	    RECT 82.6000 70.0000 106.0000 70.6000 ;
	    RECT 112.0000 70.0000 112.8000 70.6000 ;
	    RECT 82.6000 69.8000 83.6000 70.0000 ;
	    RECT 82.8000 69.6000 83.6000 69.8000 ;
	    RECT 87.6000 69.6000 88.4000 70.0000 ;
	    RECT 105.2000 69.4000 106.0000 70.0000 ;
	    RECT 71.6000 68.3000 72.4000 68.4000 ;
	    RECT 73.2000 68.3000 74.0000 68.4000 ;
	    RECT 71.6000 67.7000 74.0000 68.3000 ;
	    RECT 71.6000 67.6000 72.4000 67.7000 ;
	    RECT 73.2000 67.6000 74.0000 67.7000 ;
	    RECT 74.8000 67.6000 77.4000 68.4000 ;
	    RECT 79.6000 68.2000 80.4000 68.4000 ;
	    RECT 78.8000 67.6000 80.4000 68.2000 ;
	    RECT 81.2000 68.2000 90.0000 69.0000 ;
	    RECT 90.6000 68.6000 92.6000 69.4000 ;
	    RECT 96.4000 68.6000 99.6000 69.4000 ;
	    RECT 71.6000 64.2000 72.2000 67.6000 ;
	    RECT 73.2000 66.3000 74.0000 66.4000 ;
	    RECT 75.0000 66.3000 75.6000 67.6000 ;
	    RECT 78.8000 67.2000 79.6000 67.6000 ;
	    RECT 73.2000 65.7000 75.6000 66.3000 ;
	    RECT 76.6000 66.2000 80.2000 66.6000 ;
	    RECT 73.2000 64.8000 74.0000 65.7000 ;
	    RECT 71.6000 62.2000 72.4000 64.2000 ;
	    RECT 74.8000 62.2000 75.6000 65.7000 ;
	    RECT 76.4000 66.0000 80.4000 66.2000 ;
	    RECT 76.4000 62.2000 77.2000 66.0000 ;
	    RECT 79.6000 62.2000 80.4000 66.0000 ;
	    RECT 81.2000 62.2000 82.0000 68.2000 ;
	    RECT 83.6000 66.8000 86.6000 67.6000 ;
	    RECT 85.8000 66.2000 86.6000 66.8000 ;
	    RECT 91.8000 66.2000 92.6000 68.6000 ;
	    RECT 94.0000 66.8000 94.8000 68.4000 ;
	    RECT 99.2000 67.8000 100.0000 68.0000 ;
	    RECT 95.6000 67.2000 100.0000 67.8000 ;
	    RECT 95.6000 67.0000 96.4000 67.2000 ;
	    RECT 102.0000 66.4000 102.8000 69.2000 ;
	    RECT 107.8000 68.6000 111.6000 69.4000 ;
	    RECT 107.8000 67.4000 108.6000 68.6000 ;
	    RECT 112.2000 68.0000 112.8000 70.0000 ;
	    RECT 95.6000 66.2000 96.4000 66.4000 ;
	    RECT 85.8000 65.4000 88.4000 66.2000 ;
	    RECT 91.8000 65.6000 96.4000 66.2000 ;
	    RECT 97.2000 65.6000 98.8000 66.4000 ;
	    RECT 101.8000 65.6000 102.8000 66.4000 ;
	    RECT 106.8000 66.8000 108.6000 67.4000 ;
	    RECT 111.6000 67.4000 112.8000 68.0000 ;
	    RECT 106.8000 66.2000 107.6000 66.8000 ;
	    RECT 87.6000 62.2000 88.4000 65.4000 ;
	    RECT 105.2000 65.4000 107.6000 66.2000 ;
	    RECT 89.2000 62.2000 90.0000 65.0000 ;
	    RECT 90.8000 62.2000 91.6000 65.0000 ;
	    RECT 92.4000 62.2000 93.2000 65.0000 ;
	    RECT 95.6000 62.2000 96.4000 65.0000 ;
	    RECT 98.8000 62.2000 99.6000 65.0000 ;
	    RECT 100.4000 62.2000 101.2000 65.0000 ;
	    RECT 102.0000 62.2000 102.8000 65.0000 ;
	    RECT 103.6000 62.2000 104.4000 65.0000 ;
	    RECT 105.2000 62.2000 106.0000 65.4000 ;
	    RECT 111.6000 62.2000 112.4000 67.4000 ;
	    RECT 113.4000 66.8000 114.2000 71.2000 ;
	    RECT 113.2000 66.0000 114.2000 66.8000 ;
	    RECT 113.2000 62.2000 114.0000 66.0000 ;
	    RECT 116.4000 64.8000 117.2000 66.4000 ;
	    RECT 118.0000 62.2000 118.8000 79.8000 ;
	    RECT 119.6000 62.2000 120.4000 79.8000 ;
	    RECT 122.8000 72.4000 123.6000 79.8000 ;
	    RECT 126.0000 79.2000 130.0000 79.8000 ;
	    RECT 126.0000 72.4000 126.8000 79.2000 ;
	    RECT 122.8000 71.8000 126.8000 72.4000 ;
	    RECT 127.6000 71.8000 128.4000 78.6000 ;
	    RECT 129.2000 71.8000 130.0000 79.2000 ;
	    RECT 130.8000 73.8000 131.6000 79.8000 ;
	    RECT 131.0000 73.2000 131.6000 73.8000 ;
	    RECT 134.0000 79.2000 138.0000 79.8000 ;
	    RECT 134.0000 73.8000 134.8000 79.2000 ;
	    RECT 135.6000 73.8000 136.4000 78.6000 ;
	    RECT 137.2000 74.0000 138.0000 79.2000 ;
	    RECT 139.0000 79.2000 142.6000 79.8000 ;
	    RECT 139.0000 79.0000 139.6000 79.2000 ;
	    RECT 134.0000 73.2000 134.6000 73.8000 ;
	    RECT 131.0000 72.6000 134.6000 73.2000 ;
	    RECT 135.8000 73.4000 136.4000 73.8000 ;
	    RECT 138.8000 73.4000 139.6000 79.0000 ;
	    RECT 142.0000 79.0000 142.6000 79.2000 ;
	    RECT 135.8000 73.0000 139.6000 73.4000 ;
	    RECT 140.4000 73.0000 141.2000 78.6000 ;
	    RECT 142.0000 73.0000 142.8000 79.0000 ;
	    RECT 150.0000 76.4000 150.8000 79.8000 ;
	    RECT 149.8000 75.8000 150.8000 76.4000 ;
	    RECT 149.8000 75.2000 150.4000 75.8000 ;
	    RECT 153.2000 75.2000 154.0000 79.8000 ;
	    RECT 156.4000 77.0000 157.2000 79.8000 ;
	    RECT 158.0000 77.0000 158.8000 79.8000 ;
	    RECT 148.4000 74.6000 150.4000 75.2000 ;
	    RECT 135.8000 72.8000 139.4000 73.0000 ;
	    RECT 140.4000 72.4000 141.0000 73.0000 ;
	    RECT 140.4000 72.2000 141.2000 72.4000 ;
	    RECT 127.6000 71.2000 128.2000 71.8000 ;
	    RECT 137.8000 71.6000 141.2000 72.2000 ;
	    RECT 123.6000 70.4000 124.4000 70.8000 ;
	    RECT 126.2000 70.6000 128.2000 71.2000 ;
	    RECT 126.2000 70.4000 126.8000 70.6000 ;
	    RECT 122.8000 69.8000 124.4000 70.4000 ;
	    RECT 122.8000 69.6000 123.6000 69.8000 ;
	    RECT 126.0000 69.6000 126.8000 70.4000 ;
	    RECT 129.2000 70.3000 130.0000 71.2000 ;
	    RECT 135.6000 70.3000 137.2000 70.4000 ;
	    RECT 129.2000 69.7000 137.2000 70.3000 ;
	    RECT 129.2000 69.6000 130.0000 69.7000 ;
	    RECT 135.6000 69.6000 137.2000 69.7000 ;
	    RECT 124.4000 67.6000 125.2000 69.2000 ;
	    RECT 121.2000 64.8000 122.0000 66.4000 ;
	    RECT 126.2000 66.2000 126.8000 69.6000 ;
	    RECT 127.4000 68.8000 128.2000 69.6000 ;
	    RECT 127.6000 68.4000 128.2000 68.8000 ;
	    RECT 127.6000 67.6000 128.4000 68.4000 ;
	    RECT 132.4000 68.3000 133.2000 68.4000 ;
	    RECT 134.0000 68.3000 135.6000 68.4000 ;
	    RECT 132.4000 67.7000 135.6000 68.3000 ;
	    RECT 132.4000 67.6000 133.2000 67.7000 ;
	    RECT 134.0000 67.6000 135.6000 67.7000 ;
	    RECT 132.4000 66.3000 134.2000 66.4000 ;
	    RECT 135.6000 66.3000 136.4000 66.4000 ;
	    RECT 125.8000 64.4000 127.4000 66.2000 ;
	    RECT 132.4000 65.7000 136.4000 66.3000 ;
	    RECT 132.4000 65.6000 134.2000 65.7000 ;
	    RECT 135.6000 65.6000 136.4000 65.7000 ;
	    RECT 137.8000 65.0000 138.4000 71.6000 ;
	    RECT 134.4000 64.4000 138.4000 65.0000 ;
	    RECT 125.8000 63.6000 128.4000 64.4000 ;
	    RECT 134.0000 63.6000 135.0000 64.4000 ;
	    RECT 137.2000 64.2000 138.4000 64.4000 ;
	    RECT 148.4000 69.0000 149.2000 74.6000 ;
	    RECT 151.0000 74.4000 155.2000 75.2000 ;
	    RECT 159.6000 75.0000 160.4000 79.8000 ;
	    RECT 162.8000 75.0000 163.6000 79.8000 ;
	    RECT 151.0000 74.0000 151.6000 74.4000 ;
	    RECT 150.0000 73.2000 151.6000 74.0000 ;
	    RECT 154.6000 73.8000 160.4000 74.4000 ;
	    RECT 152.6000 73.2000 154.0000 73.8000 ;
	    RECT 152.6000 73.0000 158.8000 73.2000 ;
	    RECT 153.4000 72.6000 158.8000 73.0000 ;
	    RECT 158.0000 72.4000 158.8000 72.6000 ;
	    RECT 159.8000 73.0000 160.4000 73.8000 ;
	    RECT 161.0000 73.6000 163.6000 74.4000 ;
	    RECT 166.0000 73.6000 166.8000 79.8000 ;
	    RECT 167.6000 77.0000 168.4000 79.8000 ;
	    RECT 169.2000 77.0000 170.0000 79.8000 ;
	    RECT 170.8000 77.0000 171.6000 79.8000 ;
	    RECT 169.2000 74.4000 173.4000 75.2000 ;
	    RECT 174.0000 74.4000 174.8000 79.8000 ;
	    RECT 177.2000 75.2000 178.0000 79.8000 ;
	    RECT 177.2000 74.6000 179.8000 75.2000 ;
	    RECT 174.0000 73.6000 176.6000 74.4000 ;
	    RECT 167.6000 73.0000 168.4000 73.2000 ;
	    RECT 159.8000 72.4000 168.4000 73.0000 ;
	    RECT 170.8000 73.0000 171.6000 73.2000 ;
	    RECT 179.2000 73.0000 179.8000 74.6000 ;
	    RECT 170.8000 72.4000 179.8000 73.0000 ;
	    RECT 179.2000 70.6000 179.8000 72.4000 ;
	    RECT 180.4000 72.0000 181.2000 79.8000 ;
	    RECT 186.2000 72.4000 187.0000 79.8000 ;
	    RECT 192.6000 78.4000 193.4000 79.8000 ;
	    RECT 191.6000 77.6000 193.4000 78.4000 ;
	    RECT 187.6000 73.6000 188.4000 74.4000 ;
	    RECT 187.8000 72.4000 188.4000 73.6000 ;
	    RECT 192.6000 72.4000 193.4000 77.6000 ;
	    RECT 194.0000 73.6000 194.8000 74.4000 ;
	    RECT 194.2000 72.4000 194.8000 73.6000 ;
	    RECT 180.4000 71.2000 181.4000 72.0000 ;
	    RECT 185.2000 71.6000 187.2000 72.4000 ;
	    RECT 187.8000 71.8000 189.2000 72.4000 ;
	    RECT 192.6000 71.8000 193.6000 72.4000 ;
	    RECT 194.2000 71.8000 195.6000 72.4000 ;
	    RECT 196.4000 71.8000 197.2000 79.8000 ;
	    RECT 198.0000 72.4000 198.8000 79.8000 ;
	    RECT 201.2000 72.4000 202.0000 79.8000 ;
	    RECT 205.0000 74.4000 205.8000 79.8000 ;
	    RECT 210.8000 75.6000 211.6000 79.8000 ;
	    RECT 214.0000 75.8000 214.8000 79.8000 ;
	    RECT 214.0000 75.6000 214.6000 75.8000 ;
	    RECT 211.0000 75.0000 214.6000 75.6000 ;
	    RECT 203.6000 73.6000 204.4000 74.4000 ;
	    RECT 205.0000 73.6000 206.8000 74.4000 ;
	    RECT 203.6000 72.4000 204.2000 73.6000 ;
	    RECT 205.0000 72.4000 205.8000 73.6000 ;
	    RECT 212.4000 72.8000 213.2000 74.4000 ;
	    RECT 214.0000 72.4000 214.6000 75.0000 ;
	    RECT 218.2000 74.4000 219.0000 79.8000 ;
	    RECT 217.2000 73.6000 219.0000 74.4000 ;
	    RECT 218.2000 72.4000 219.0000 73.6000 ;
	    RECT 222.6000 78.4000 223.4000 79.8000 ;
	    RECT 222.6000 77.6000 224.4000 78.4000 ;
	    RECT 222.6000 72.6000 223.4000 77.6000 ;
	    RECT 198.0000 71.8000 202.0000 72.4000 ;
	    RECT 202.8000 71.8000 204.2000 72.4000 ;
	    RECT 204.8000 71.8000 205.8000 72.4000 ;
	    RECT 188.4000 71.6000 189.2000 71.8000 ;
	    RECT 149.8000 70.0000 173.2000 70.6000 ;
	    RECT 179.2000 70.0000 180.0000 70.6000 ;
	    RECT 149.8000 69.8000 150.6000 70.0000 ;
	    RECT 151.6000 69.6000 152.4000 70.0000 ;
	    RECT 154.8000 69.6000 155.6000 70.0000 ;
	    RECT 161.2000 69.6000 162.0000 70.0000 ;
	    RECT 172.4000 69.4000 173.2000 70.0000 ;
	    RECT 148.4000 68.2000 157.2000 69.0000 ;
	    RECT 157.8000 68.6000 159.8000 69.4000 ;
	    RECT 163.6000 68.6000 166.8000 69.4000 ;
	    RECT 125.8000 62.2000 127.4000 63.6000 ;
	    RECT 134.0000 62.2000 134.8000 63.6000 ;
	    RECT 137.2000 62.2000 138.0000 64.2000 ;
	    RECT 148.4000 62.2000 149.2000 68.2000 ;
	    RECT 150.8000 66.8000 153.8000 67.6000 ;
	    RECT 153.0000 66.2000 153.8000 66.8000 ;
	    RECT 159.0000 66.2000 159.8000 68.6000 ;
	    RECT 161.2000 66.8000 162.0000 68.4000 ;
	    RECT 166.4000 67.8000 167.2000 68.0000 ;
	    RECT 162.8000 67.2000 167.2000 67.8000 ;
	    RECT 162.8000 67.0000 163.6000 67.2000 ;
	    RECT 169.2000 66.4000 170.0000 69.2000 ;
	    RECT 175.0000 68.6000 178.8000 69.4000 ;
	    RECT 175.0000 67.4000 175.8000 68.6000 ;
	    RECT 179.4000 68.0000 180.0000 70.0000 ;
	    RECT 162.8000 66.2000 163.6000 66.4000 ;
	    RECT 153.0000 65.4000 155.6000 66.2000 ;
	    RECT 159.0000 65.6000 163.6000 66.2000 ;
	    RECT 164.4000 65.6000 166.0000 66.4000 ;
	    RECT 169.0000 65.6000 170.0000 66.4000 ;
	    RECT 174.0000 66.8000 175.8000 67.4000 ;
	    RECT 178.8000 67.4000 180.0000 68.0000 ;
	    RECT 174.0000 66.2000 174.8000 66.8000 ;
	    RECT 154.8000 62.2000 155.6000 65.4000 ;
	    RECT 172.4000 65.4000 174.8000 66.2000 ;
	    RECT 156.4000 62.2000 157.2000 65.0000 ;
	    RECT 158.0000 62.2000 158.8000 65.0000 ;
	    RECT 159.6000 62.2000 160.4000 65.0000 ;
	    RECT 162.8000 62.2000 163.6000 65.0000 ;
	    RECT 166.0000 62.2000 166.8000 65.0000 ;
	    RECT 167.6000 62.2000 168.4000 65.0000 ;
	    RECT 169.2000 62.2000 170.0000 65.0000 ;
	    RECT 170.8000 62.2000 171.6000 65.0000 ;
	    RECT 172.4000 62.2000 173.2000 65.4000 ;
	    RECT 178.8000 62.2000 179.6000 67.4000 ;
	    RECT 180.6000 66.8000 181.4000 71.2000 ;
	    RECT 185.2000 68.8000 186.0000 70.4000 ;
	    RECT 186.6000 68.4000 187.2000 71.6000 ;
	    RECT 191.6000 68.8000 192.4000 70.4000 ;
	    RECT 193.0000 68.4000 193.6000 71.8000 ;
	    RECT 194.8000 71.6000 195.6000 71.8000 ;
	    RECT 196.6000 70.4000 197.2000 71.8000 ;
	    RECT 202.8000 71.6000 203.6000 71.8000 ;
	    RECT 200.4000 70.4000 201.2000 70.8000 ;
	    RECT 196.4000 69.8000 198.8000 70.4000 ;
	    RECT 200.4000 69.8000 202.0000 70.4000 ;
	    RECT 196.4000 69.6000 197.2000 69.8000 ;
	    RECT 198.0000 69.6000 198.8000 69.8000 ;
	    RECT 201.2000 69.6000 202.0000 69.8000 ;
	    RECT 183.6000 68.2000 184.4000 68.4000 ;
	    RECT 183.6000 67.6000 185.2000 68.2000 ;
	    RECT 186.6000 67.6000 189.2000 68.4000 ;
	    RECT 190.0000 68.2000 190.8000 68.4000 ;
	    RECT 190.0000 67.6000 191.6000 68.2000 ;
	    RECT 193.0000 67.6000 195.6000 68.4000 ;
	    RECT 184.4000 67.2000 185.2000 67.6000 ;
	    RECT 180.4000 66.0000 181.4000 66.8000 ;
	    RECT 183.8000 66.2000 187.4000 66.6000 ;
	    RECT 188.4000 66.2000 189.0000 67.6000 ;
	    RECT 190.8000 67.2000 191.6000 67.6000 ;
	    RECT 190.2000 66.2000 193.8000 66.6000 ;
	    RECT 194.8000 66.2000 195.4000 67.6000 ;
	    RECT 183.6000 66.0000 187.6000 66.2000 ;
	    RECT 180.4000 62.2000 181.2000 66.0000 ;
	    RECT 183.6000 62.2000 184.4000 66.0000 ;
	    RECT 186.8000 62.2000 187.6000 66.0000 ;
	    RECT 188.4000 62.2000 189.2000 66.2000 ;
	    RECT 190.0000 66.0000 194.0000 66.2000 ;
	    RECT 190.0000 62.2000 190.8000 66.0000 ;
	    RECT 193.2000 62.2000 194.0000 66.0000 ;
	    RECT 194.8000 62.2000 195.6000 66.2000 ;
	    RECT 196.4000 65.6000 197.2000 66.4000 ;
	    RECT 198.2000 66.2000 198.8000 69.6000 ;
	    RECT 204.8000 68.4000 205.4000 71.8000 ;
	    RECT 209.2000 70.8000 210.0000 72.4000 ;
	    RECT 214.0000 71.6000 214.8000 72.4000 ;
	    RECT 218.2000 71.8000 219.2000 72.4000 ;
	    RECT 222.6000 71.8000 224.4000 72.6000 ;
	    RECT 206.0000 68.8000 206.8000 70.4000 ;
	    RECT 210.8000 69.6000 212.4000 70.4000 ;
	    RECT 214.0000 68.4000 214.6000 71.6000 ;
	    RECT 217.2000 68.8000 218.0000 70.4000 ;
	    RECT 202.8000 67.6000 205.4000 68.4000 ;
	    RECT 213.0000 68.2000 214.6000 68.4000 ;
	    RECT 212.8000 67.8000 214.6000 68.2000 ;
	    RECT 218.6000 68.4000 219.2000 71.8000 ;
	    RECT 223.6000 68.4000 224.2000 71.8000 ;
	    RECT 203.0000 66.2000 203.6000 67.6000 ;
	    RECT 204.6000 66.2000 208.2000 66.6000 ;
	    RECT 196.6000 64.8000 197.4000 65.6000 ;
	    RECT 198.0000 62.2000 198.8000 66.2000 ;
	    RECT 202.8000 62.2000 203.6000 66.2000 ;
	    RECT 204.4000 66.0000 208.4000 66.2000 ;
	    RECT 204.4000 62.2000 205.2000 66.0000 ;
	    RECT 207.6000 62.2000 208.4000 66.0000 ;
	    RECT 212.8000 62.2000 213.6000 67.8000 ;
	    RECT 218.6000 67.6000 221.2000 68.4000 ;
	    RECT 223.6000 67.6000 224.4000 68.4000 ;
	    RECT 215.8000 66.2000 219.4000 66.6000 ;
	    RECT 220.4000 66.2000 221.0000 67.6000 ;
	    RECT 215.6000 66.0000 219.6000 66.2000 ;
	    RECT 215.6000 62.2000 216.4000 66.0000 ;
	    RECT 218.8000 62.2000 219.6000 66.0000 ;
	    RECT 220.4000 62.2000 221.2000 66.2000 ;
	    RECT 223.6000 64.2000 224.2000 67.6000 ;
	    RECT 223.6000 62.2000 224.4000 64.2000 ;
	    RECT 4.4000 55.2000 5.2000 59.8000 ;
	    RECT 9.2000 55.2000 10.0000 59.8000 ;
	    RECT 14.6000 56.0000 15.4000 59.0000 ;
	    RECT 18.8000 57.0000 19.6000 59.0000 ;
	    RECT 3.0000 54.6000 5.2000 55.2000 ;
	    RECT 7.8000 54.6000 10.0000 55.2000 ;
	    RECT 13.8000 55.4000 15.4000 56.0000 ;
	    RECT 13.8000 55.0000 14.6000 55.4000 ;
	    RECT 3.0000 51.6000 3.6000 54.6000 ;
	    RECT 4.4000 51.6000 5.2000 53.2000 ;
	    RECT 7.8000 51.6000 8.4000 54.6000 ;
	    RECT 13.8000 54.4000 14.4000 55.0000 ;
	    RECT 19.0000 54.8000 19.6000 57.0000 ;
	    RECT 12.4000 53.6000 14.4000 54.4000 ;
	    RECT 15.4000 54.2000 19.6000 54.8000 ;
	    RECT 20.4000 54.3000 21.2000 59.8000 ;
	    RECT 22.0000 55.6000 22.8000 57.2000 ;
	    RECT 26.8000 55.8000 27.6000 59.8000 ;
	    RECT 28.2000 56.4000 29.0000 57.2000 ;
	    RECT 25.2000 54.3000 26.0000 54.4000 ;
	    RECT 15.4000 53.8000 16.4000 54.2000 ;
	    RECT 9.2000 51.6000 10.0000 53.2000 ;
	    RECT 2.4000 50.8000 3.6000 51.6000 ;
	    RECT 7.2000 50.8000 8.4000 51.6000 ;
	    RECT 12.4000 50.8000 13.2000 52.4000 ;
	    RECT 3.0000 50.2000 3.6000 50.8000 ;
	    RECT 7.8000 50.2000 8.4000 50.8000 ;
	    RECT 3.0000 49.6000 5.2000 50.2000 ;
	    RECT 7.8000 49.6000 10.0000 50.2000 ;
	    RECT 4.4000 42.2000 5.2000 49.6000 ;
	    RECT 9.2000 42.2000 10.0000 49.6000 ;
	    RECT 13.8000 49.8000 14.4000 53.6000 ;
	    RECT 15.0000 53.0000 16.4000 53.8000 ;
	    RECT 20.4000 53.7000 26.0000 54.3000 ;
	    RECT 15.8000 51.0000 16.4000 53.0000 ;
	    RECT 17.2000 51.6000 18.0000 53.2000 ;
	    RECT 18.8000 51.6000 19.6000 53.2000 ;
	    RECT 15.8000 50.4000 19.6000 51.0000 ;
	    RECT 13.8000 49.2000 15.4000 49.8000 ;
	    RECT 14.6000 44.4000 15.4000 49.2000 ;
	    RECT 19.0000 47.0000 19.6000 50.4000 ;
	    RECT 14.0000 43.6000 15.4000 44.4000 ;
	    RECT 14.6000 42.2000 15.4000 43.6000 ;
	    RECT 18.8000 43.0000 19.6000 47.0000 ;
	    RECT 20.4000 42.2000 21.2000 53.7000 ;
	    RECT 25.2000 52.8000 26.0000 53.7000 ;
	    RECT 23.6000 52.2000 24.4000 52.4000 ;
	    RECT 26.8000 52.2000 27.4000 55.8000 ;
	    RECT 28.4000 55.6000 29.2000 56.4000 ;
	    RECT 33.2000 55.8000 34.0000 59.8000 ;
	    RECT 34.6000 56.4000 35.4000 57.2000 ;
	    RECT 31.6000 52.8000 32.4000 54.4000 ;
	    RECT 28.4000 52.2000 29.2000 52.4000 ;
	    RECT 23.6000 51.6000 25.2000 52.2000 ;
	    RECT 26.8000 51.6000 29.2000 52.2000 ;
	    RECT 30.0000 52.2000 30.8000 52.4000 ;
	    RECT 33.2000 52.2000 33.8000 55.8000 ;
	    RECT 34.8000 55.6000 35.6000 56.4000 ;
	    RECT 34.8000 52.2000 35.6000 52.4000 ;
	    RECT 30.0000 51.6000 31.6000 52.2000 ;
	    RECT 33.2000 51.6000 35.6000 52.2000 ;
	    RECT 24.4000 51.2000 25.2000 51.6000 ;
	    RECT 28.4000 50.2000 29.0000 51.6000 ;
	    RECT 30.8000 51.2000 31.6000 51.6000 ;
	    RECT 34.8000 50.2000 35.4000 51.6000 ;
	    RECT 23.6000 49.6000 27.6000 50.2000 ;
	    RECT 23.6000 42.2000 24.4000 49.6000 ;
	    RECT 26.8000 42.2000 27.6000 49.6000 ;
	    RECT 28.4000 42.2000 29.2000 50.2000 ;
	    RECT 30.0000 49.6000 34.0000 50.2000 ;
	    RECT 30.0000 42.2000 30.8000 49.6000 ;
	    RECT 33.2000 42.2000 34.0000 49.6000 ;
	    RECT 34.8000 42.2000 35.6000 50.2000 ;
	    RECT 36.4000 42.2000 37.2000 59.8000 ;
	    RECT 38.0000 55.6000 38.8000 57.2000 ;
	    RECT 39.6000 55.8000 40.4000 59.8000 ;
	    RECT 44.0000 58.4000 45.6000 59.8000 ;
	    RECT 44.0000 57.6000 46.8000 58.4000 ;
	    RECT 44.0000 56.2000 45.6000 57.6000 ;
	    RECT 38.1000 54.4000 38.7000 55.6000 ;
	    RECT 39.6000 55.2000 42.0000 55.8000 ;
	    RECT 41.2000 55.0000 42.0000 55.2000 ;
	    RECT 42.6000 54.8000 43.4000 55.6000 ;
	    RECT 42.6000 54.4000 43.2000 54.8000 ;
	    RECT 38.0000 54.3000 38.8000 54.4000 ;
	    RECT 39.6000 54.3000 41.2000 54.4000 ;
	    RECT 38.0000 53.7000 41.2000 54.3000 ;
	    RECT 38.0000 53.6000 38.8000 53.7000 ;
	    RECT 39.6000 53.6000 41.2000 53.7000 ;
	    RECT 42.4000 53.6000 43.2000 54.4000 ;
	    RECT 44.0000 52.8000 44.6000 56.2000 ;
	    RECT 49.2000 55.8000 50.0000 59.8000 ;
	    RECT 45.2000 55.4000 46.8000 55.6000 ;
	    RECT 45.2000 54.8000 47.2000 55.4000 ;
	    RECT 47.8000 55.2000 50.0000 55.8000 ;
	    RECT 50.8000 57.0000 51.6000 59.0000 ;
	    RECT 47.8000 55.0000 48.6000 55.2000 ;
	    RECT 46.6000 54.4000 47.2000 54.8000 ;
	    RECT 50.8000 54.8000 51.4000 57.0000 ;
	    RECT 55.0000 56.0000 55.8000 59.0000 ;
	    RECT 55.0000 55.4000 56.6000 56.0000 ;
	    RECT 55.8000 55.0000 56.6000 55.4000 ;
	    RECT 45.2000 53.4000 46.0000 54.2000 ;
	    RECT 46.6000 53.8000 50.0000 54.4000 ;
	    RECT 50.8000 54.2000 55.0000 54.8000 ;
	    RECT 48.4000 53.6000 50.0000 53.8000 ;
	    RECT 54.0000 53.8000 55.0000 54.2000 ;
	    RECT 56.0000 54.4000 56.6000 55.0000 ;
	    RECT 43.6000 52.4000 44.6000 52.8000 ;
	    RECT 42.8000 52.2000 44.6000 52.4000 ;
	    RECT 45.4000 52.8000 46.0000 53.4000 ;
	    RECT 45.4000 52.2000 48.0000 52.8000 ;
	    RECT 42.8000 51.6000 44.2000 52.2000 ;
	    RECT 47.2000 52.0000 48.0000 52.2000 ;
	    RECT 50.8000 51.6000 51.6000 53.2000 ;
	    RECT 52.4000 51.6000 53.2000 53.2000 ;
	    RECT 54.0000 53.0000 55.4000 53.8000 ;
	    RECT 56.0000 53.6000 58.0000 54.4000 ;
	    RECT 43.6000 50.2000 44.2000 51.6000 ;
	    RECT 45.0000 51.4000 45.8000 51.6000 ;
	    RECT 45.0000 50.8000 48.4000 51.4000 ;
	    RECT 54.0000 51.0000 54.6000 53.0000 ;
	    RECT 47.8000 50.2000 48.4000 50.8000 ;
	    RECT 50.8000 50.4000 54.6000 51.0000 ;
	    RECT 39.6000 49.6000 42.0000 50.2000 ;
	    RECT 43.6000 49.6000 45.6000 50.2000 ;
	    RECT 39.6000 42.2000 40.4000 49.6000 ;
	    RECT 41.2000 49.4000 42.0000 49.6000 ;
	    RECT 44.0000 42.2000 45.6000 49.6000 ;
	    RECT 47.8000 49.6000 50.0000 50.2000 ;
	    RECT 47.8000 49.4000 48.6000 49.6000 ;
	    RECT 49.2000 42.2000 50.0000 49.6000 ;
	    RECT 50.8000 47.0000 51.4000 50.4000 ;
	    RECT 56.0000 49.8000 56.6000 53.6000 ;
	    RECT 60.4000 52.4000 61.2000 59.8000 ;
	    RECT 63.6000 55.2000 64.4000 59.8000 ;
	    RECT 62.2000 54.6000 64.4000 55.2000 ;
	    RECT 57.2000 50.8000 58.0000 52.4000 ;
	    RECT 55.0000 49.2000 56.6000 49.8000 ;
	    RECT 60.4000 50.2000 61.0000 52.4000 ;
	    RECT 62.2000 51.6000 62.8000 54.6000 ;
	    RECT 63.6000 52.3000 64.4000 53.2000 ;
	    RECT 68.4000 52.3000 69.2000 52.4000 ;
	    RECT 63.6000 51.7000 69.2000 52.3000 ;
	    RECT 63.6000 51.6000 64.4000 51.7000 ;
	    RECT 68.4000 51.6000 69.2000 51.7000 ;
	    RECT 61.6000 50.8000 62.8000 51.6000 ;
	    RECT 62.2000 50.2000 62.8000 50.8000 ;
	    RECT 50.8000 43.0000 51.6000 47.0000 ;
	    RECT 55.0000 44.4000 55.8000 49.2000 ;
	    RECT 55.0000 43.6000 56.4000 44.4000 ;
	    RECT 55.0000 42.2000 55.8000 43.6000 ;
	    RECT 60.4000 42.2000 61.2000 50.2000 ;
	    RECT 62.2000 49.6000 64.4000 50.2000 ;
	    RECT 63.6000 42.2000 64.4000 49.6000 ;
	    RECT 70.0000 42.2000 70.8000 59.8000 ;
	    RECT 71.6000 55.6000 72.4000 57.2000 ;
	    RECT 74.8000 55.2000 75.6000 59.8000 ;
	    RECT 78.0000 55.2000 78.8000 59.8000 ;
	    RECT 81.2000 55.2000 82.0000 59.8000 ;
	    RECT 84.4000 55.2000 85.2000 59.8000 ;
	    RECT 73.2000 54.4000 75.6000 55.2000 ;
	    RECT 76.6000 54.4000 78.8000 55.2000 ;
	    RECT 79.8000 54.4000 82.0000 55.2000 ;
	    RECT 83.4000 54.4000 85.2000 55.2000 ;
	    RECT 89.2000 55.2000 90.0000 59.8000 ;
	    RECT 92.4000 55.2000 93.2000 59.8000 ;
	    RECT 95.6000 55.2000 96.4000 59.8000 ;
	    RECT 98.8000 55.2000 99.6000 59.8000 ;
	    RECT 103.6000 57.6000 104.4000 59.8000 ;
	    RECT 102.0000 55.6000 102.8000 57.2000 ;
	    RECT 89.2000 54.4000 91.0000 55.2000 ;
	    RECT 92.4000 54.4000 94.6000 55.2000 ;
	    RECT 95.6000 54.4000 97.8000 55.2000 ;
	    RECT 98.8000 54.4000 101.2000 55.2000 ;
	    RECT 103.8000 54.4000 104.4000 57.6000 ;
	    RECT 107.4000 56.4000 108.2000 59.8000 ;
	    RECT 107.4000 55.8000 109.2000 56.4000 ;
	    RECT 73.2000 51.6000 74.0000 54.4000 ;
	    RECT 76.6000 53.8000 77.4000 54.4000 ;
	    RECT 79.8000 53.8000 80.6000 54.4000 ;
	    RECT 83.4000 53.8000 84.2000 54.4000 ;
	    RECT 74.8000 53.0000 77.4000 53.8000 ;
	    RECT 78.2000 53.0000 80.6000 53.8000 ;
	    RECT 81.6000 53.0000 84.2000 53.8000 ;
	    RECT 76.6000 51.6000 77.4000 53.0000 ;
	    RECT 79.8000 51.6000 80.6000 53.0000 ;
	    RECT 83.4000 51.6000 84.2000 53.0000 ;
	    RECT 90.2000 53.8000 91.0000 54.4000 ;
	    RECT 93.8000 53.8000 94.6000 54.4000 ;
	    RECT 97.0000 53.8000 97.8000 54.4000 ;
	    RECT 90.2000 53.0000 92.8000 53.8000 ;
	    RECT 93.8000 53.0000 96.2000 53.8000 ;
	    RECT 97.0000 53.0000 99.6000 53.8000 ;
	    RECT 90.2000 51.6000 91.0000 53.0000 ;
	    RECT 93.8000 51.6000 94.6000 53.0000 ;
	    RECT 97.0000 51.6000 97.8000 53.0000 ;
	    RECT 100.4000 51.6000 101.2000 54.4000 ;
	    RECT 103.6000 53.6000 104.4000 54.4000 ;
	    RECT 73.2000 50.8000 75.6000 51.6000 ;
	    RECT 76.6000 50.8000 78.8000 51.6000 ;
	    RECT 79.8000 50.8000 82.0000 51.6000 ;
	    RECT 83.4000 50.8000 85.2000 51.6000 ;
	    RECT 74.8000 42.2000 75.6000 50.8000 ;
	    RECT 78.0000 42.2000 78.8000 50.8000 ;
	    RECT 81.2000 42.2000 82.0000 50.8000 ;
	    RECT 84.4000 42.2000 85.2000 50.8000 ;
	    RECT 89.2000 50.8000 91.0000 51.6000 ;
	    RECT 92.4000 50.8000 94.6000 51.6000 ;
	    RECT 95.6000 50.8000 97.8000 51.6000 ;
	    RECT 98.8000 50.8000 101.2000 51.6000 ;
	    RECT 89.2000 42.2000 90.0000 50.8000 ;
	    RECT 92.4000 42.2000 93.2000 50.8000 ;
	    RECT 95.6000 42.2000 96.4000 50.8000 ;
	    RECT 98.8000 42.2000 99.6000 50.8000 ;
	    RECT 103.8000 50.2000 104.4000 53.6000 ;
	    RECT 105.2000 52.3000 106.0000 52.4000 ;
	    RECT 108.4000 52.3000 109.2000 55.8000 ;
	    RECT 110.0000 53.6000 110.8000 55.2000 ;
	    RECT 115.2000 54.2000 116.0000 59.8000 ;
	    RECT 119.2000 54.2000 120.0000 59.8000 ;
	    RECT 126.0000 56.0000 126.8000 59.8000 ;
	    RECT 115.2000 53.8000 117.0000 54.2000 ;
	    RECT 115.4000 53.6000 117.0000 53.8000 ;
	    RECT 105.2000 51.7000 109.2000 52.3000 ;
	    RECT 110.1000 52.3000 110.7000 53.6000 ;
	    RECT 110.1000 51.7000 112.4000 52.3000 ;
	    RECT 105.2000 50.8000 106.0000 51.7000 ;
	    RECT 103.6000 49.4000 105.4000 50.2000 ;
	    RECT 104.6000 44.4000 105.4000 49.4000 ;
	    RECT 106.8000 48.8000 107.6000 50.4000 ;
	    RECT 103.6000 43.6000 105.4000 44.4000 ;
	    RECT 104.6000 42.2000 105.4000 43.6000 ;
	    RECT 108.4000 42.2000 109.2000 51.7000 ;
	    RECT 111.6000 49.6000 112.4000 51.7000 ;
	    RECT 113.2000 51.6000 114.8000 52.4000 ;
	    RECT 116.4000 50.4000 117.0000 53.6000 ;
	    RECT 118.2000 53.8000 120.0000 54.2000 ;
	    RECT 125.8000 55.2000 126.8000 56.0000 ;
	    RECT 118.2000 53.6000 119.8000 53.8000 ;
	    RECT 118.2000 50.4000 118.8000 53.6000 ;
	    RECT 120.4000 51.6000 122.0000 52.4000 ;
	    RECT 116.4000 49.6000 117.2000 50.4000 ;
	    RECT 118.0000 49.6000 118.8000 50.4000 ;
	    RECT 122.8000 49.6000 123.6000 51.2000 ;
	    RECT 125.8000 50.8000 126.6000 55.2000 ;
	    RECT 127.6000 54.6000 128.4000 59.8000 ;
	    RECT 134.0000 56.6000 134.8000 59.8000 ;
	    RECT 135.6000 57.0000 136.4000 59.8000 ;
	    RECT 137.2000 57.0000 138.0000 59.8000 ;
	    RECT 138.8000 57.0000 139.6000 59.8000 ;
	    RECT 140.4000 57.0000 141.2000 59.8000 ;
	    RECT 143.6000 57.0000 144.4000 59.8000 ;
	    RECT 146.8000 57.0000 147.6000 59.8000 ;
	    RECT 148.4000 57.0000 149.2000 59.8000 ;
	    RECT 150.0000 57.0000 150.8000 59.8000 ;
	    RECT 132.4000 55.8000 134.8000 56.6000 ;
	    RECT 151.6000 56.6000 152.4000 59.8000 ;
	    RECT 132.4000 55.2000 133.2000 55.8000 ;
	    RECT 127.2000 54.0000 128.4000 54.6000 ;
	    RECT 131.4000 54.6000 133.2000 55.2000 ;
	    RECT 137.2000 55.6000 138.2000 56.4000 ;
	    RECT 141.2000 55.6000 142.8000 56.4000 ;
	    RECT 143.6000 55.8000 148.2000 56.4000 ;
	    RECT 151.6000 55.8000 154.2000 56.6000 ;
	    RECT 143.6000 55.6000 144.4000 55.8000 ;
	    RECT 127.2000 52.0000 127.8000 54.0000 ;
	    RECT 131.4000 53.4000 132.2000 54.6000 ;
	    RECT 128.4000 52.6000 132.2000 53.4000 ;
	    RECT 137.2000 52.8000 138.0000 55.6000 ;
	    RECT 143.6000 54.8000 144.4000 55.0000 ;
	    RECT 140.0000 54.2000 144.4000 54.8000 ;
	    RECT 140.0000 54.0000 140.8000 54.2000 ;
	    RECT 145.2000 53.6000 146.0000 55.2000 ;
	    RECT 147.4000 53.4000 148.2000 55.8000 ;
	    RECT 153.4000 55.2000 154.2000 55.8000 ;
	    RECT 153.4000 54.4000 156.4000 55.2000 ;
	    RECT 158.0000 53.8000 158.8000 59.8000 ;
	    RECT 164.4000 56.0000 165.2000 59.8000 ;
	    RECT 167.6000 56.0000 168.4000 59.8000 ;
	    RECT 164.4000 55.8000 168.4000 56.0000 ;
	    RECT 169.2000 55.8000 170.0000 59.8000 ;
	    RECT 170.8000 55.8000 171.6000 59.8000 ;
	    RECT 175.0000 58.4000 175.8000 59.8000 ;
	    RECT 175.0000 57.6000 176.4000 58.4000 ;
	    RECT 175.0000 56.8000 175.8000 57.6000 ;
	    RECT 175.0000 55.8000 176.4000 56.8000 ;
	    RECT 177.2000 55.8000 178.0000 59.8000 ;
	    RECT 178.8000 56.0000 179.6000 59.8000 ;
	    RECT 182.0000 56.0000 182.8000 59.8000 ;
	    RECT 178.8000 55.8000 182.8000 56.0000 ;
	    RECT 185.2000 57.8000 186.0000 59.8000 ;
	    RECT 164.6000 55.4000 168.2000 55.8000 ;
	    RECT 165.2000 54.4000 166.0000 54.8000 ;
	    RECT 169.2000 54.4000 169.8000 55.8000 ;
	    RECT 171.0000 55.6000 171.6000 55.8000 ;
	    RECT 171.0000 55.2000 172.8000 55.6000 ;
	    RECT 171.0000 55.0000 175.2000 55.2000 ;
	    RECT 172.2000 54.6000 175.2000 55.0000 ;
	    RECT 174.4000 54.4000 175.2000 54.6000 ;
	    RECT 140.4000 52.6000 143.6000 53.4000 ;
	    RECT 147.4000 52.6000 149.4000 53.4000 ;
	    RECT 150.0000 53.0000 158.8000 53.8000 ;
	    RECT 164.4000 53.8000 166.0000 54.4000 ;
	    RECT 164.4000 53.6000 165.2000 53.8000 ;
	    RECT 167.4000 53.6000 170.0000 54.4000 ;
	    RECT 134.0000 52.0000 134.8000 52.6000 ;
	    RECT 151.6000 52.0000 152.4000 52.4000 ;
	    RECT 156.6000 52.0000 157.4000 52.2000 ;
	    RECT 127.2000 51.4000 128.0000 52.0000 ;
	    RECT 134.0000 51.4000 157.4000 52.0000 ;
	    RECT 125.8000 50.0000 126.8000 50.8000 ;
	    RECT 114.8000 47.6000 115.6000 49.2000 ;
	    RECT 116.4000 47.0000 117.0000 49.6000 ;
	    RECT 113.4000 46.4000 117.0000 47.0000 ;
	    RECT 113.4000 46.2000 114.0000 46.4000 ;
	    RECT 113.2000 42.2000 114.0000 46.2000 ;
	    RECT 116.4000 46.2000 117.0000 46.4000 ;
	    RECT 118.2000 47.0000 118.8000 49.6000 ;
	    RECT 119.6000 47.6000 120.4000 49.2000 ;
	    RECT 118.2000 46.4000 121.8000 47.0000 ;
	    RECT 118.2000 46.2000 118.8000 46.4000 ;
	    RECT 116.4000 42.2000 117.2000 46.2000 ;
	    RECT 118.0000 42.2000 118.8000 46.2000 ;
	    RECT 121.2000 42.2000 122.0000 46.4000 ;
	    RECT 126.0000 42.2000 126.8000 50.0000 ;
	    RECT 127.4000 49.6000 128.0000 51.4000 ;
	    RECT 127.4000 49.0000 136.4000 49.6000 ;
	    RECT 127.4000 47.4000 128.0000 49.0000 ;
	    RECT 135.6000 48.8000 136.4000 49.0000 ;
	    RECT 138.8000 49.0000 147.4000 49.6000 ;
	    RECT 138.8000 48.8000 139.6000 49.0000 ;
	    RECT 130.6000 47.6000 133.2000 48.4000 ;
	    RECT 127.4000 46.8000 130.0000 47.4000 ;
	    RECT 129.2000 42.2000 130.0000 46.8000 ;
	    RECT 132.4000 42.2000 133.2000 47.6000 ;
	    RECT 133.8000 46.8000 138.0000 47.6000 ;
	    RECT 135.6000 42.2000 136.4000 45.0000 ;
	    RECT 137.2000 42.2000 138.0000 45.0000 ;
	    RECT 138.8000 42.2000 139.6000 45.0000 ;
	    RECT 140.4000 42.2000 141.2000 48.4000 ;
	    RECT 143.6000 47.6000 146.2000 48.4000 ;
	    RECT 146.8000 48.2000 147.4000 49.0000 ;
	    RECT 148.4000 49.4000 149.2000 49.6000 ;
	    RECT 148.4000 49.0000 153.8000 49.4000 ;
	    RECT 148.4000 48.8000 154.6000 49.0000 ;
	    RECT 153.2000 48.2000 154.6000 48.8000 ;
	    RECT 146.8000 47.6000 152.6000 48.2000 ;
	    RECT 155.6000 48.0000 157.2000 48.8000 ;
	    RECT 155.6000 47.6000 156.2000 48.0000 ;
	    RECT 143.6000 42.2000 144.4000 47.0000 ;
	    RECT 146.8000 42.2000 147.6000 47.0000 ;
	    RECT 152.0000 46.8000 156.2000 47.6000 ;
	    RECT 158.0000 47.4000 158.8000 53.0000 ;
	    RECT 166.0000 51.6000 166.8000 53.2000 ;
	    RECT 167.4000 50.2000 168.0000 53.6000 ;
	    RECT 170.8000 52.8000 171.6000 54.4000 ;
	    RECT 172.8000 53.8000 173.6000 54.0000 ;
	    RECT 172.6000 53.2000 173.6000 53.8000 ;
	    RECT 172.6000 52.4000 173.2000 53.2000 ;
	    RECT 172.4000 51.6000 173.2000 52.4000 ;
	    RECT 174.4000 51.0000 175.0000 54.4000 ;
	    RECT 175.8000 52.4000 176.4000 55.8000 ;
	    RECT 177.4000 54.4000 178.0000 55.8000 ;
	    RECT 179.0000 55.4000 182.6000 55.8000 ;
	    RECT 181.2000 54.4000 182.0000 54.8000 ;
	    RECT 185.2000 54.4000 185.8000 57.8000 ;
	    RECT 186.8000 55.6000 187.6000 57.2000 ;
	    RECT 188.4000 55.8000 189.2000 59.8000 ;
	    RECT 192.8000 58.4000 194.4000 59.8000 ;
	    RECT 191.6000 57.6000 194.4000 58.4000 ;
	    RECT 192.8000 56.2000 194.4000 57.6000 ;
	    RECT 188.4000 55.2000 191.0000 55.8000 ;
	    RECT 190.2000 55.0000 191.0000 55.2000 ;
	    RECT 191.6000 54.8000 193.2000 55.6000 ;
	    RECT 177.2000 53.6000 179.8000 54.4000 ;
	    RECT 181.2000 53.8000 182.8000 54.4000 ;
	    RECT 182.0000 53.6000 182.8000 53.8000 ;
	    RECT 185.2000 53.6000 186.0000 54.4000 ;
	    RECT 188.4000 54.2000 190.0000 54.4000 ;
	    RECT 193.8000 54.2000 194.4000 56.2000 ;
	    RECT 198.0000 55.8000 198.8000 59.8000 ;
	    RECT 199.6000 55.8000 200.4000 59.8000 ;
	    RECT 201.2000 56.0000 202.0000 59.8000 ;
	    RECT 204.4000 56.0000 205.2000 59.8000 ;
	    RECT 201.2000 55.8000 205.2000 56.0000 ;
	    RECT 195.0000 54.8000 195.8000 55.6000 ;
	    RECT 196.4000 55.2000 198.8000 55.8000 ;
	    RECT 196.4000 55.0000 197.2000 55.2000 ;
	    RECT 188.4000 54.0000 190.6000 54.2000 ;
	    RECT 188.4000 53.6000 192.8000 54.0000 ;
	    RECT 175.6000 51.6000 176.4000 52.4000 ;
	    RECT 172.6000 50.4000 175.0000 51.0000 ;
	    RECT 169.2000 50.2000 170.0000 50.4000 ;
	    RECT 156.8000 46.8000 158.8000 47.4000 ;
	    RECT 167.0000 49.6000 168.0000 50.2000 ;
	    RECT 168.6000 49.6000 170.0000 50.2000 ;
	    RECT 148.4000 42.2000 149.2000 45.0000 ;
	    RECT 150.0000 42.2000 150.8000 45.0000 ;
	    RECT 153.2000 42.2000 154.0000 46.8000 ;
	    RECT 156.8000 46.2000 157.4000 46.8000 ;
	    RECT 156.4000 45.6000 157.4000 46.2000 ;
	    RECT 156.4000 42.2000 157.2000 45.6000 ;
	    RECT 167.0000 42.2000 167.8000 49.6000 ;
	    RECT 168.6000 48.4000 169.2000 49.6000 ;
	    RECT 168.4000 47.6000 169.2000 48.4000 ;
	    RECT 172.6000 46.2000 173.2000 50.4000 ;
	    RECT 175.8000 50.2000 176.4000 51.6000 ;
	    RECT 172.4000 42.2000 173.2000 46.2000 ;
	    RECT 175.6000 42.2000 176.4000 50.2000 ;
	    RECT 177.2000 50.2000 178.0000 50.4000 ;
	    RECT 179.2000 50.2000 179.8000 53.6000 ;
	    RECT 180.4000 51.6000 181.2000 53.2000 ;
	    RECT 182.1000 52.3000 182.7000 53.6000 ;
	    RECT 183.6000 52.3000 184.4000 52.4000 ;
	    RECT 182.1000 51.7000 184.4000 52.3000 ;
	    RECT 183.6000 50.8000 184.4000 51.7000 ;
	    RECT 185.2000 50.2000 185.8000 53.6000 ;
	    RECT 190.0000 53.4000 192.8000 53.6000 ;
	    RECT 192.0000 53.2000 192.8000 53.4000 ;
	    RECT 193.4000 53.6000 194.4000 54.2000 ;
	    RECT 195.2000 54.4000 195.8000 54.8000 ;
	    RECT 199.8000 54.4000 200.4000 55.8000 ;
	    RECT 201.4000 55.4000 205.0000 55.8000 ;
	    RECT 206.0000 55.2000 206.8000 59.8000 ;
	    RECT 210.8000 55.6000 211.6000 57.2000 ;
	    RECT 203.6000 54.4000 204.4000 54.8000 ;
	    RECT 206.0000 54.6000 208.2000 55.2000 ;
	    RECT 195.2000 53.6000 196.0000 54.4000 ;
	    RECT 197.2000 53.6000 198.8000 54.4000 ;
	    RECT 199.6000 53.6000 202.2000 54.4000 ;
	    RECT 203.6000 53.8000 205.2000 54.4000 ;
	    RECT 204.4000 53.6000 205.2000 53.8000 ;
	    RECT 193.4000 52.4000 194.0000 53.6000 ;
	    RECT 190.6000 52.2000 191.4000 52.4000 ;
	    RECT 190.6000 51.6000 192.2000 52.2000 ;
	    RECT 193.2000 51.6000 194.0000 52.4000 ;
	    RECT 194.8000 52.3000 195.6000 52.4000 ;
	    RECT 201.6000 52.3000 202.2000 53.6000 ;
	    RECT 194.8000 51.7000 202.2000 52.3000 ;
	    RECT 194.8000 51.6000 195.6000 51.7000 ;
	    RECT 191.4000 51.4000 192.2000 51.6000 ;
	    RECT 193.4000 50.2000 194.0000 51.6000 ;
	    RECT 199.6000 50.2000 200.4000 50.4000 ;
	    RECT 201.6000 50.2000 202.2000 51.7000 ;
	    RECT 202.8000 51.6000 203.6000 53.2000 ;
	    RECT 204.4000 52.3000 205.2000 52.4000 ;
	    RECT 206.0000 52.3000 206.8000 53.2000 ;
	    RECT 204.4000 51.7000 206.8000 52.3000 ;
	    RECT 204.4000 51.6000 205.2000 51.7000 ;
	    RECT 206.0000 51.6000 206.8000 51.7000 ;
	    RECT 207.6000 51.6000 208.2000 54.6000 ;
	    RECT 207.6000 50.8000 208.8000 51.6000 ;
	    RECT 207.6000 50.2000 208.2000 50.8000 ;
	    RECT 177.2000 49.6000 178.6000 50.2000 ;
	    RECT 179.2000 49.6000 180.2000 50.2000 ;
	    RECT 178.0000 48.4000 178.6000 49.6000 ;
	    RECT 178.0000 47.6000 178.8000 48.4000 ;
	    RECT 179.4000 42.2000 180.2000 49.6000 ;
	    RECT 184.2000 49.4000 186.0000 50.2000 ;
	    RECT 188.4000 49.6000 191.0000 50.2000 ;
	    RECT 184.2000 48.4000 185.0000 49.4000 ;
	    RECT 183.6000 47.6000 185.0000 48.4000 ;
	    RECT 184.2000 42.2000 185.0000 47.6000 ;
	    RECT 188.4000 42.2000 189.2000 49.6000 ;
	    RECT 190.2000 49.4000 191.0000 49.6000 ;
	    RECT 192.8000 42.2000 194.4000 50.2000 ;
	    RECT 196.4000 49.6000 198.8000 50.2000 ;
	    RECT 199.6000 49.6000 201.0000 50.2000 ;
	    RECT 201.6000 49.6000 202.6000 50.2000 ;
	    RECT 196.4000 49.4000 197.2000 49.6000 ;
	    RECT 198.0000 42.2000 198.8000 49.6000 ;
	    RECT 200.4000 48.4000 201.0000 49.6000 ;
	    RECT 200.4000 47.6000 201.2000 48.4000 ;
	    RECT 201.8000 42.2000 202.6000 49.6000 ;
	    RECT 206.0000 49.6000 208.2000 50.2000 ;
	    RECT 206.0000 42.2000 206.8000 49.6000 ;
	    RECT 212.4000 42.2000 213.2000 59.8000 ;
	    RECT 215.6000 57.8000 216.4000 59.8000 ;
	    RECT 219.4000 58.4000 220.2000 59.8000 ;
	    RECT 215.8000 54.4000 216.4000 57.8000 ;
	    RECT 218.8000 57.6000 220.2000 58.4000 ;
	    RECT 219.4000 56.4000 220.2000 57.6000 ;
	    RECT 217.2000 56.3000 218.0000 56.4000 ;
	    RECT 219.4000 56.3000 221.2000 56.4000 ;
	    RECT 217.2000 55.7000 221.2000 56.3000 ;
	    RECT 217.2000 55.6000 218.0000 55.7000 ;
	    RECT 214.0000 54.3000 214.8000 54.4000 ;
	    RECT 215.6000 54.3000 216.4000 54.4000 ;
	    RECT 214.0000 53.7000 216.4000 54.3000 ;
	    RECT 214.0000 53.6000 214.8000 53.7000 ;
	    RECT 215.6000 53.6000 216.4000 53.7000 ;
	    RECT 215.8000 50.2000 216.4000 53.6000 ;
	    RECT 215.6000 49.4000 217.4000 50.2000 ;
	    RECT 216.6000 42.2000 217.4000 49.4000 ;
	    RECT 220.4000 42.2000 221.2000 55.7000 ;
	    RECT 1.2000 24.8000 2.0000 26.4000 ;
	    RECT 2.8000 22.2000 3.6000 39.8000 ;
	    RECT 6.0000 32.0000 6.8000 39.8000 ;
	    RECT 9.2000 35.2000 10.0000 39.8000 ;
	    RECT 5.8000 31.2000 6.8000 32.0000 ;
	    RECT 7.4000 34.6000 10.0000 35.2000 ;
	    RECT 7.4000 33.0000 8.0000 34.6000 ;
	    RECT 12.4000 34.4000 13.2000 39.8000 ;
	    RECT 15.6000 37.0000 16.4000 39.8000 ;
	    RECT 17.2000 37.0000 18.0000 39.8000 ;
	    RECT 18.8000 37.0000 19.6000 39.8000 ;
	    RECT 13.8000 34.4000 18.0000 35.2000 ;
	    RECT 10.6000 33.6000 13.2000 34.4000 ;
	    RECT 20.4000 33.6000 21.2000 39.8000 ;
	    RECT 23.6000 35.0000 24.4000 39.8000 ;
	    RECT 26.8000 35.0000 27.6000 39.8000 ;
	    RECT 28.4000 37.0000 29.2000 39.8000 ;
	    RECT 30.0000 37.0000 30.8000 39.8000 ;
	    RECT 33.2000 35.2000 34.0000 39.8000 ;
	    RECT 36.4000 36.4000 37.2000 39.8000 ;
	    RECT 41.2000 36.4000 42.0000 39.8000 ;
	    RECT 36.4000 35.8000 37.4000 36.4000 ;
	    RECT 36.8000 35.2000 37.4000 35.8000 ;
	    RECT 41.0000 35.8000 42.0000 36.4000 ;
	    RECT 41.0000 35.2000 41.6000 35.8000 ;
	    RECT 44.4000 35.2000 45.2000 39.8000 ;
	    RECT 47.6000 37.0000 48.4000 39.8000 ;
	    RECT 49.2000 37.0000 50.0000 39.8000 ;
	    RECT 32.0000 34.4000 36.2000 35.2000 ;
	    RECT 36.8000 34.6000 38.8000 35.2000 ;
	    RECT 23.6000 33.6000 26.2000 34.4000 ;
	    RECT 26.8000 33.8000 32.6000 34.4000 ;
	    RECT 35.6000 34.0000 36.2000 34.4000 ;
	    RECT 15.6000 33.0000 16.4000 33.2000 ;
	    RECT 7.4000 32.4000 16.4000 33.0000 ;
	    RECT 18.8000 33.0000 19.6000 33.2000 ;
	    RECT 26.8000 33.0000 27.4000 33.8000 ;
	    RECT 33.2000 33.2000 34.6000 33.8000 ;
	    RECT 35.6000 33.2000 37.2000 34.0000 ;
	    RECT 18.8000 32.4000 27.4000 33.0000 ;
	    RECT 28.4000 33.0000 34.6000 33.2000 ;
	    RECT 28.4000 32.6000 33.8000 33.0000 ;
	    RECT 28.4000 32.4000 29.2000 32.6000 ;
	    RECT 5.8000 26.8000 6.6000 31.2000 ;
	    RECT 7.4000 30.6000 8.0000 32.4000 ;
	    RECT 7.2000 30.0000 8.0000 30.6000 ;
	    RECT 14.0000 30.0000 37.4000 30.6000 ;
	    RECT 7.2000 28.0000 7.8000 30.0000 ;
	    RECT 14.0000 29.4000 14.8000 30.0000 ;
	    RECT 31.6000 29.6000 32.4000 30.0000 ;
	    RECT 33.2000 29.6000 34.0000 30.0000 ;
	    RECT 34.8000 29.6000 35.6000 30.0000 ;
	    RECT 36.6000 29.8000 37.4000 30.0000 ;
	    RECT 8.4000 28.6000 12.2000 29.4000 ;
	    RECT 7.2000 27.4000 8.4000 28.0000 ;
	    RECT 5.8000 26.0000 6.8000 26.8000 ;
	    RECT 6.0000 22.2000 6.8000 26.0000 ;
	    RECT 7.6000 22.2000 8.4000 27.4000 ;
	    RECT 11.4000 27.4000 12.2000 28.6000 ;
	    RECT 11.4000 26.8000 13.2000 27.4000 ;
	    RECT 12.4000 26.2000 13.2000 26.8000 ;
	    RECT 17.2000 26.4000 18.0000 29.2000 ;
	    RECT 20.4000 28.6000 23.6000 29.4000 ;
	    RECT 27.4000 28.6000 29.4000 29.4000 ;
	    RECT 38.0000 29.0000 38.8000 34.6000 ;
	    RECT 20.0000 27.8000 20.8000 28.0000 ;
	    RECT 20.0000 27.2000 24.4000 27.8000 ;
	    RECT 23.6000 27.0000 24.4000 27.2000 ;
	    RECT 25.2000 26.8000 26.0000 28.4000 ;
	    RECT 12.4000 25.4000 14.8000 26.2000 ;
	    RECT 17.2000 25.6000 18.2000 26.4000 ;
	    RECT 21.2000 25.6000 22.8000 26.4000 ;
	    RECT 23.6000 26.2000 24.4000 26.4000 ;
	    RECT 27.4000 26.2000 28.2000 28.6000 ;
	    RECT 30.0000 28.2000 38.8000 29.0000 ;
	    RECT 33.4000 26.8000 36.4000 27.6000 ;
	    RECT 33.4000 26.2000 34.2000 26.8000 ;
	    RECT 23.6000 25.6000 28.2000 26.2000 ;
	    RECT 14.0000 22.2000 14.8000 25.4000 ;
	    RECT 31.6000 25.4000 34.2000 26.2000 ;
	    RECT 15.6000 22.2000 16.4000 25.0000 ;
	    RECT 17.2000 22.2000 18.0000 25.0000 ;
	    RECT 18.8000 22.2000 19.6000 25.0000 ;
	    RECT 20.4000 22.2000 21.2000 25.0000 ;
	    RECT 23.6000 22.2000 24.4000 25.0000 ;
	    RECT 26.8000 22.2000 27.6000 25.0000 ;
	    RECT 28.4000 22.2000 29.2000 25.0000 ;
	    RECT 30.0000 22.2000 30.8000 25.0000 ;
	    RECT 31.6000 22.2000 32.4000 25.4000 ;
	    RECT 38.0000 22.2000 38.8000 28.2000 ;
	    RECT 39.6000 34.6000 41.6000 35.2000 ;
	    RECT 39.6000 29.0000 40.4000 34.6000 ;
	    RECT 42.2000 34.4000 46.4000 35.2000 ;
	    RECT 50.8000 35.0000 51.6000 39.8000 ;
	    RECT 54.0000 35.0000 54.8000 39.8000 ;
	    RECT 42.2000 34.0000 42.8000 34.4000 ;
	    RECT 41.2000 33.2000 42.8000 34.0000 ;
	    RECT 45.8000 33.8000 51.6000 34.4000 ;
	    RECT 43.8000 33.2000 45.2000 33.8000 ;
	    RECT 43.8000 33.0000 50.0000 33.2000 ;
	    RECT 44.6000 32.6000 50.0000 33.0000 ;
	    RECT 49.2000 32.4000 50.0000 32.6000 ;
	    RECT 51.0000 33.0000 51.6000 33.8000 ;
	    RECT 52.2000 33.6000 54.8000 34.4000 ;
	    RECT 57.2000 33.6000 58.0000 39.8000 ;
	    RECT 58.8000 37.0000 59.6000 39.8000 ;
	    RECT 60.4000 37.0000 61.2000 39.8000 ;
	    RECT 62.0000 37.0000 62.8000 39.8000 ;
	    RECT 60.4000 34.4000 64.6000 35.2000 ;
	    RECT 65.2000 34.4000 66.0000 39.8000 ;
	    RECT 68.4000 35.2000 69.2000 39.8000 ;
	    RECT 68.4000 34.6000 71.0000 35.2000 ;
	    RECT 65.2000 33.6000 67.8000 34.4000 ;
	    RECT 58.8000 33.0000 59.6000 33.2000 ;
	    RECT 51.0000 32.4000 59.6000 33.0000 ;
	    RECT 62.0000 33.0000 62.8000 33.2000 ;
	    RECT 70.4000 33.0000 71.0000 34.6000 ;
	    RECT 62.0000 32.4000 71.0000 33.0000 ;
	    RECT 70.4000 30.6000 71.0000 32.4000 ;
	    RECT 71.6000 32.0000 72.4000 39.8000 ;
	    RECT 71.6000 31.2000 72.6000 32.0000 ;
	    RECT 41.0000 30.0000 64.4000 30.6000 ;
	    RECT 70.4000 30.0000 71.2000 30.6000 ;
	    RECT 41.0000 29.8000 41.8000 30.0000 ;
	    RECT 44.4000 29.6000 45.2000 30.0000 ;
	    RECT 46.0000 29.6000 46.8000 30.0000 ;
	    RECT 63.6000 29.4000 64.4000 30.0000 ;
	    RECT 39.6000 28.2000 48.4000 29.0000 ;
	    RECT 49.0000 28.6000 51.0000 29.4000 ;
	    RECT 54.8000 28.6000 58.0000 29.4000 ;
	    RECT 39.6000 22.2000 40.4000 28.2000 ;
	    RECT 42.0000 26.8000 45.0000 27.6000 ;
	    RECT 44.2000 26.2000 45.0000 26.8000 ;
	    RECT 50.2000 26.2000 51.0000 28.6000 ;
	    RECT 52.4000 26.8000 53.2000 28.4000 ;
	    RECT 57.6000 27.8000 58.4000 28.0000 ;
	    RECT 54.0000 27.2000 58.4000 27.8000 ;
	    RECT 54.0000 27.0000 54.8000 27.2000 ;
	    RECT 60.4000 26.4000 61.2000 29.2000 ;
	    RECT 66.2000 28.6000 70.0000 29.4000 ;
	    RECT 66.2000 27.4000 67.0000 28.6000 ;
	    RECT 70.6000 28.0000 71.2000 30.0000 ;
	    RECT 54.0000 26.2000 54.8000 26.4000 ;
	    RECT 44.2000 25.4000 46.8000 26.2000 ;
	    RECT 50.2000 25.6000 54.8000 26.2000 ;
	    RECT 55.6000 25.6000 57.2000 26.4000 ;
	    RECT 60.2000 25.6000 61.2000 26.4000 ;
	    RECT 65.2000 26.8000 67.0000 27.4000 ;
	    RECT 70.0000 27.4000 71.2000 28.0000 ;
	    RECT 65.2000 26.2000 66.0000 26.8000 ;
	    RECT 46.0000 22.2000 46.8000 25.4000 ;
	    RECT 63.6000 25.4000 66.0000 26.2000 ;
	    RECT 47.6000 22.2000 48.4000 25.0000 ;
	    RECT 49.2000 22.2000 50.0000 25.0000 ;
	    RECT 50.8000 22.2000 51.6000 25.0000 ;
	    RECT 54.0000 22.2000 54.8000 25.0000 ;
	    RECT 57.2000 22.2000 58.0000 25.0000 ;
	    RECT 58.8000 22.2000 59.6000 25.0000 ;
	    RECT 60.4000 22.2000 61.2000 25.0000 ;
	    RECT 62.0000 22.2000 62.8000 25.0000 ;
	    RECT 63.6000 22.2000 64.4000 25.4000 ;
	    RECT 70.0000 22.2000 70.8000 27.4000 ;
	    RECT 71.8000 26.8000 72.6000 31.2000 ;
	    RECT 79.6000 26.8000 80.4000 28.4000 ;
	    RECT 71.6000 26.0000 72.6000 26.8000 ;
	    RECT 81.2000 26.2000 82.0000 39.8000 ;
	    RECT 84.4000 33.6000 86.0000 34.4000 ;
	    RECT 82.8000 31.6000 83.6000 33.2000 ;
	    RECT 85.2000 32.4000 85.8000 33.6000 ;
	    RECT 86.6000 32.4000 87.4000 39.8000 ;
	    RECT 84.4000 31.8000 85.8000 32.4000 ;
	    RECT 86.4000 31.8000 87.4000 32.4000 ;
	    RECT 93.4000 32.4000 94.2000 39.8000 ;
	    RECT 94.8000 33.6000 95.6000 34.4000 ;
	    RECT 95.0000 32.4000 95.6000 33.6000 ;
	    RECT 93.4000 31.8000 94.4000 32.4000 ;
	    RECT 95.0000 32.3000 96.4000 32.4000 ;
	    RECT 97.2000 32.3000 98.0000 32.4000 ;
	    RECT 95.0000 31.8000 98.0000 32.3000 ;
	    RECT 84.4000 31.6000 85.2000 31.8000 ;
	    RECT 82.9000 30.3000 83.5000 31.6000 ;
	    RECT 86.4000 30.3000 87.0000 31.8000 ;
	    RECT 82.9000 29.7000 87.0000 30.3000 ;
	    RECT 86.4000 28.4000 87.0000 29.7000 ;
	    RECT 87.6000 30.3000 88.4000 30.4000 ;
	    RECT 92.4000 30.3000 93.2000 30.4000 ;
	    RECT 87.6000 29.7000 93.2000 30.3000 ;
	    RECT 87.6000 28.8000 88.4000 29.7000 ;
	    RECT 92.4000 28.8000 93.2000 29.7000 ;
	    RECT 93.8000 28.4000 94.4000 31.8000 ;
	    RECT 95.6000 31.7000 98.0000 31.8000 ;
	    RECT 95.6000 31.6000 96.4000 31.7000 ;
	    RECT 97.2000 31.6000 98.0000 31.7000 ;
	    RECT 84.4000 27.6000 87.0000 28.4000 ;
	    RECT 89.2000 28.2000 90.0000 28.4000 ;
	    RECT 88.4000 27.6000 90.0000 28.2000 ;
	    RECT 90.8000 28.2000 91.6000 28.4000 ;
	    RECT 90.8000 27.6000 92.4000 28.2000 ;
	    RECT 93.8000 27.6000 96.4000 28.4000 ;
	    RECT 84.6000 26.2000 85.2000 27.6000 ;
	    RECT 88.4000 27.2000 89.2000 27.6000 ;
	    RECT 91.6000 27.2000 92.4000 27.6000 ;
	    RECT 86.2000 26.2000 89.8000 26.6000 ;
	    RECT 91.0000 26.2000 94.6000 26.6000 ;
	    RECT 95.6000 26.2000 96.2000 27.6000 ;
	    RECT 71.6000 22.2000 72.4000 26.0000 ;
	    RECT 81.2000 25.6000 83.0000 26.2000 ;
	    RECT 82.2000 22.2000 83.0000 25.6000 ;
	    RECT 84.4000 22.2000 85.2000 26.2000 ;
	    RECT 86.0000 26.0000 90.0000 26.2000 ;
	    RECT 86.0000 22.2000 86.8000 26.0000 ;
	    RECT 89.2000 22.2000 90.0000 26.0000 ;
	    RECT 90.8000 26.0000 94.8000 26.2000 ;
	    RECT 90.8000 22.2000 91.6000 26.0000 ;
	    RECT 94.0000 22.2000 94.8000 26.0000 ;
	    RECT 95.6000 22.2000 96.4000 26.2000 ;
	    RECT 97.2000 24.8000 98.0000 26.4000 ;
	    RECT 98.8000 22.2000 99.6000 39.8000 ;
	    RECT 102.0000 35.8000 102.8000 39.8000 ;
	    RECT 102.2000 35.6000 102.8000 35.8000 ;
	    RECT 105.2000 35.6000 106.0000 39.8000 ;
	    RECT 106.8000 35.8000 107.6000 39.8000 ;
	    RECT 107.0000 35.6000 107.6000 35.8000 ;
	    RECT 110.0000 35.8000 110.8000 39.8000 ;
	    RECT 110.0000 35.6000 110.6000 35.8000 ;
	    RECT 102.2000 35.0000 105.8000 35.6000 ;
	    RECT 103.6000 32.8000 104.4000 34.4000 ;
	    RECT 105.2000 32.4000 105.8000 35.0000 ;
	    RECT 107.0000 35.0000 110.6000 35.6000 ;
	    RECT 107.0000 32.4000 107.6000 35.0000 ;
	    RECT 108.4000 32.8000 109.2000 34.4000 ;
	    RECT 100.4000 30.8000 101.2000 32.4000 ;
	    RECT 105.2000 31.6000 106.0000 32.4000 ;
	    RECT 106.8000 31.6000 107.6000 32.4000 ;
	    RECT 102.0000 29.6000 103.6000 30.4000 ;
	    RECT 105.2000 28.4000 105.8000 31.6000 ;
	    RECT 104.2000 28.2000 105.8000 28.4000 ;
	    RECT 104.0000 27.8000 105.8000 28.2000 ;
	    RECT 107.0000 28.4000 107.6000 31.6000 ;
	    RECT 111.6000 30.8000 112.4000 32.4000 ;
	    RECT 113.2000 31.8000 114.0000 39.8000 ;
	    RECT 116.4000 35.8000 117.2000 39.8000 ;
	    RECT 113.2000 30.4000 113.8000 31.8000 ;
	    RECT 116.4000 31.6000 117.0000 35.8000 ;
	    RECT 122.2000 32.6000 123.0000 39.8000 ;
	    RECT 121.2000 31.8000 123.0000 32.6000 ;
	    RECT 126.0000 32.0000 126.8000 39.8000 ;
	    RECT 129.2000 35.2000 130.0000 39.8000 ;
	    RECT 114.6000 31.0000 117.0000 31.6000 ;
	    RECT 109.2000 29.6000 110.8000 30.4000 ;
	    RECT 113.2000 29.6000 114.0000 30.4000 ;
	    RECT 107.0000 28.2000 108.6000 28.4000 ;
	    RECT 107.0000 27.8000 108.8000 28.2000 ;
	    RECT 104.0000 22.2000 104.8000 27.8000 ;
	    RECT 108.0000 26.3000 108.8000 27.8000 ;
	    RECT 110.0000 26.3000 110.8000 26.4000 ;
	    RECT 108.0000 25.7000 110.8000 26.3000 ;
	    RECT 108.0000 22.2000 108.8000 25.7000 ;
	    RECT 110.0000 25.6000 110.8000 25.7000 ;
	    RECT 113.2000 26.2000 113.8000 29.6000 ;
	    RECT 114.6000 27.6000 115.2000 31.0000 ;
	    RECT 116.4000 29.6000 117.2000 30.4000 ;
	    RECT 119.6000 30.3000 120.4000 30.4000 ;
	    RECT 121.4000 30.3000 122.0000 31.8000 ;
	    RECT 125.8000 31.2000 126.8000 32.0000 ;
	    RECT 127.4000 34.6000 130.0000 35.2000 ;
	    RECT 127.4000 33.0000 128.0000 34.6000 ;
	    RECT 132.4000 34.4000 133.2000 39.8000 ;
	    RECT 135.6000 37.0000 136.4000 39.8000 ;
	    RECT 137.2000 37.0000 138.0000 39.8000 ;
	    RECT 138.8000 37.0000 139.6000 39.8000 ;
	    RECT 133.8000 34.4000 138.0000 35.2000 ;
	    RECT 130.6000 33.6000 133.2000 34.4000 ;
	    RECT 140.4000 33.6000 141.2000 39.8000 ;
	    RECT 143.6000 35.0000 144.4000 39.8000 ;
	    RECT 146.8000 35.0000 147.6000 39.8000 ;
	    RECT 148.4000 37.0000 149.2000 39.8000 ;
	    RECT 150.0000 37.0000 150.8000 39.8000 ;
	    RECT 153.2000 35.2000 154.0000 39.8000 ;
	    RECT 156.4000 36.4000 157.2000 39.8000 ;
	    RECT 156.4000 35.8000 157.4000 36.4000 ;
	    RECT 156.8000 35.2000 157.4000 35.8000 ;
	    RECT 152.0000 34.4000 156.2000 35.2000 ;
	    RECT 156.8000 34.6000 158.8000 35.2000 ;
	    RECT 143.6000 33.6000 146.2000 34.4000 ;
	    RECT 146.8000 33.8000 152.6000 34.4000 ;
	    RECT 155.6000 34.0000 156.2000 34.4000 ;
	    RECT 135.6000 33.0000 136.4000 33.2000 ;
	    RECT 127.4000 32.4000 136.4000 33.0000 ;
	    RECT 138.8000 33.0000 139.6000 33.2000 ;
	    RECT 146.8000 33.0000 147.4000 33.8000 ;
	    RECT 153.2000 33.2000 154.6000 33.8000 ;
	    RECT 155.6000 33.2000 157.2000 34.0000 ;
	    RECT 138.8000 32.4000 147.4000 33.0000 ;
	    RECT 148.4000 33.0000 154.6000 33.2000 ;
	    RECT 148.4000 32.6000 153.8000 33.0000 ;
	    RECT 148.4000 32.4000 149.2000 32.6000 ;
	    RECT 119.6000 29.7000 122.0000 30.3000 ;
	    RECT 119.6000 29.6000 120.4000 29.7000 ;
	    RECT 116.4000 28.8000 117.0000 29.6000 ;
	    RECT 116.0000 28.2000 117.0000 28.8000 ;
	    RECT 116.0000 28.0000 116.8000 28.2000 ;
	    RECT 118.0000 27.6000 118.8000 29.2000 ;
	    RECT 121.4000 28.4000 122.0000 29.7000 ;
	    RECT 122.8000 30.3000 123.6000 31.2000 ;
	    RECT 125.8000 30.3000 126.6000 31.2000 ;
	    RECT 127.4000 30.6000 128.0000 32.4000 ;
	    RECT 122.8000 29.7000 126.6000 30.3000 ;
	    RECT 122.8000 29.6000 123.6000 29.7000 ;
	    RECT 121.2000 27.6000 122.0000 28.4000 ;
	    RECT 114.4000 27.4000 115.2000 27.6000 ;
	    RECT 114.4000 27.0000 117.4000 27.4000 ;
	    RECT 114.4000 26.8000 118.6000 27.0000 ;
	    RECT 116.8000 26.4000 118.6000 26.8000 ;
	    RECT 118.0000 26.2000 118.6000 26.4000 ;
	    RECT 113.2000 25.2000 114.6000 26.2000 ;
	    RECT 113.8000 24.4000 114.6000 25.2000 ;
	    RECT 113.2000 23.6000 114.6000 24.4000 ;
	    RECT 113.8000 22.2000 114.6000 23.6000 ;
	    RECT 118.0000 22.2000 118.8000 26.2000 ;
	    RECT 119.6000 24.8000 120.4000 26.4000 ;
	    RECT 121.4000 24.2000 122.0000 27.6000 ;
	    RECT 125.8000 26.8000 126.6000 29.7000 ;
	    RECT 127.2000 30.0000 128.0000 30.6000 ;
	    RECT 134.0000 30.0000 157.4000 30.6000 ;
	    RECT 127.2000 28.0000 127.8000 30.0000 ;
	    RECT 134.0000 29.4000 134.8000 30.0000 ;
	    RECT 151.6000 29.6000 152.4000 30.0000 ;
	    RECT 156.6000 29.8000 157.4000 30.0000 ;
	    RECT 128.4000 28.6000 132.2000 29.4000 ;
	    RECT 127.2000 27.4000 128.4000 28.0000 ;
	    RECT 125.8000 26.0000 126.8000 26.8000 ;
	    RECT 121.2000 22.2000 122.0000 24.2000 ;
	    RECT 126.0000 22.2000 126.8000 26.0000 ;
	    RECT 127.6000 22.2000 128.4000 27.4000 ;
	    RECT 131.4000 27.4000 132.2000 28.6000 ;
	    RECT 131.4000 26.8000 133.2000 27.4000 ;
	    RECT 132.4000 26.2000 133.2000 26.8000 ;
	    RECT 137.2000 26.4000 138.0000 29.2000 ;
	    RECT 140.4000 28.6000 143.6000 29.4000 ;
	    RECT 147.4000 28.6000 149.4000 29.4000 ;
	    RECT 158.0000 29.0000 158.8000 34.6000 ;
	    RECT 140.0000 27.8000 140.8000 28.0000 ;
	    RECT 140.0000 27.2000 144.4000 27.8000 ;
	    RECT 143.6000 27.0000 144.4000 27.2000 ;
	    RECT 145.2000 26.8000 146.0000 28.4000 ;
	    RECT 132.4000 25.4000 134.8000 26.2000 ;
	    RECT 137.2000 25.6000 138.2000 26.4000 ;
	    RECT 141.2000 25.6000 142.8000 26.4000 ;
	    RECT 143.6000 26.2000 144.4000 26.4000 ;
	    RECT 147.4000 26.2000 148.2000 28.6000 ;
	    RECT 150.0000 28.2000 158.8000 29.0000 ;
	    RECT 153.4000 26.8000 156.4000 27.6000 ;
	    RECT 153.4000 26.2000 154.2000 26.8000 ;
	    RECT 143.6000 25.6000 148.2000 26.2000 ;
	    RECT 134.0000 22.2000 134.8000 25.4000 ;
	    RECT 151.6000 25.4000 154.2000 26.2000 ;
	    RECT 135.6000 22.2000 136.4000 25.0000 ;
	    RECT 137.2000 22.2000 138.0000 25.0000 ;
	    RECT 138.8000 22.2000 139.6000 25.0000 ;
	    RECT 140.4000 22.2000 141.2000 25.0000 ;
	    RECT 143.6000 22.2000 144.4000 25.0000 ;
	    RECT 146.8000 22.2000 147.6000 25.0000 ;
	    RECT 148.4000 22.2000 149.2000 25.0000 ;
	    RECT 150.0000 22.2000 150.8000 25.0000 ;
	    RECT 151.6000 22.2000 152.4000 25.4000 ;
	    RECT 158.0000 22.2000 158.8000 28.2000 ;
	    RECT 166.0000 28.3000 166.8000 39.8000 ;
	    RECT 167.6000 28.3000 168.4000 28.4000 ;
	    RECT 166.0000 27.7000 168.4000 28.3000 ;
	    RECT 162.8000 26.3000 163.6000 26.4000 ;
	    RECT 164.4000 26.3000 165.2000 26.4000 ;
	    RECT 162.8000 25.7000 165.2000 26.3000 ;
	    RECT 162.8000 25.6000 163.6000 25.7000 ;
	    RECT 164.4000 24.8000 165.2000 25.7000 ;
	    RECT 166.0000 22.2000 166.8000 27.7000 ;
	    RECT 167.6000 26.8000 168.4000 27.7000 ;
	    RECT 169.2000 26.4000 170.0000 39.8000 ;
	    RECT 170.8000 31.6000 171.6000 33.2000 ;
	    RECT 173.0000 32.6000 173.8000 39.8000 ;
	    RECT 173.0000 31.8000 174.8000 32.6000 ;
	    RECT 170.9000 30.3000 171.5000 31.6000 ;
	    RECT 172.4000 30.3000 173.2000 31.2000 ;
	    RECT 170.9000 29.7000 173.2000 30.3000 ;
	    RECT 172.4000 29.6000 173.2000 29.7000 ;
	    RECT 174.0000 28.4000 174.6000 31.8000 ;
	    RECT 178.8000 30.3000 179.6000 39.8000 ;
	    RECT 183.0000 32.4000 183.8000 39.8000 ;
	    RECT 184.4000 33.6000 185.2000 34.4000 ;
	    RECT 184.6000 32.4000 185.2000 33.6000 ;
	    RECT 183.0000 31.8000 184.0000 32.4000 ;
	    RECT 184.6000 31.8000 186.0000 32.4000 ;
	    RECT 182.0000 30.3000 182.8000 30.4000 ;
	    RECT 178.8000 29.7000 182.8000 30.3000 ;
	    RECT 174.0000 28.3000 174.8000 28.4000 ;
	    RECT 177.2000 28.3000 178.0000 28.4000 ;
	    RECT 174.0000 27.7000 178.0000 28.3000 ;
	    RECT 174.0000 27.6000 174.8000 27.7000 ;
	    RECT 177.2000 27.6000 178.0000 27.7000 ;
	    RECT 169.2000 25.6000 171.6000 26.4000 ;
	    RECT 170.2000 22.2000 171.0000 25.6000 ;
	    RECT 174.0000 24.2000 174.6000 27.6000 ;
	    RECT 175.6000 24.8000 176.4000 26.4000 ;
	    RECT 177.2000 24.8000 178.0000 26.4000 ;
	    RECT 174.0000 22.2000 174.8000 24.2000 ;
	    RECT 178.8000 22.2000 179.6000 29.7000 ;
	    RECT 182.0000 28.8000 182.8000 29.7000 ;
	    RECT 183.4000 30.3000 184.0000 31.8000 ;
	    RECT 185.2000 31.6000 186.0000 31.8000 ;
	    RECT 186.8000 31.6000 187.6000 33.2000 ;
	    RECT 186.9000 30.3000 187.5000 31.6000 ;
	    RECT 183.4000 29.7000 187.5000 30.3000 ;
	    RECT 183.4000 28.4000 184.0000 29.7000 ;
	    RECT 180.4000 28.2000 181.2000 28.4000 ;
	    RECT 180.4000 27.6000 182.0000 28.2000 ;
	    RECT 183.4000 27.6000 186.0000 28.4000 ;
	    RECT 181.2000 27.2000 182.0000 27.6000 ;
	    RECT 180.6000 26.2000 184.2000 26.6000 ;
	    RECT 185.2000 26.2000 185.8000 27.6000 ;
	    RECT 188.4000 26.2000 189.2000 39.8000 ;
	    RECT 193.2000 35.6000 194.0000 39.8000 ;
	    RECT 196.4000 35.8000 197.2000 39.8000 ;
	    RECT 196.4000 35.6000 197.0000 35.8000 ;
	    RECT 193.4000 35.0000 197.0000 35.6000 ;
	    RECT 194.8000 32.8000 195.6000 34.4000 ;
	    RECT 196.4000 32.4000 197.0000 35.0000 ;
	    RECT 198.8000 33.6000 199.6000 34.4000 ;
	    RECT 198.8000 32.4000 199.4000 33.6000 ;
	    RECT 200.2000 32.4000 201.0000 39.8000 ;
	    RECT 191.6000 30.8000 192.4000 32.4000 ;
	    RECT 196.4000 31.6000 197.2000 32.4000 ;
	    RECT 198.0000 31.8000 199.4000 32.4000 ;
	    RECT 200.0000 31.8000 201.0000 32.4000 ;
	    RECT 206.0000 32.3000 206.8000 39.8000 ;
	    RECT 209.8000 38.4000 210.6000 39.8000 ;
	    RECT 209.8000 37.6000 211.6000 38.4000 ;
	    RECT 208.4000 33.6000 209.2000 34.4000 ;
	    RECT 208.4000 32.4000 209.0000 33.6000 ;
	    RECT 209.8000 32.4000 210.6000 37.6000 ;
	    RECT 215.6000 35.6000 216.4000 39.8000 ;
	    RECT 218.8000 35.8000 219.6000 39.8000 ;
	    RECT 223.0000 38.4000 223.8000 39.8000 ;
	    RECT 223.0000 37.6000 224.4000 38.4000 ;
	    RECT 218.8000 35.6000 219.4000 35.8000 ;
	    RECT 215.8000 35.0000 219.4000 35.6000 ;
	    RECT 217.2000 32.8000 218.0000 34.4000 ;
	    RECT 218.8000 32.4000 219.4000 35.0000 ;
	    RECT 223.0000 32.6000 223.8000 37.6000 ;
	    RECT 207.6000 32.3000 209.0000 32.4000 ;
	    RECT 206.0000 31.8000 209.0000 32.3000 ;
	    RECT 209.6000 31.8000 210.6000 32.4000 ;
	    RECT 198.0000 31.6000 198.8000 31.8000 ;
	    RECT 193.2000 29.6000 194.8000 30.4000 ;
	    RECT 196.4000 28.4000 197.0000 31.6000 ;
	    RECT 200.0000 28.4000 200.6000 31.8000 ;
	    RECT 206.0000 31.7000 208.4000 31.8000 ;
	    RECT 201.2000 28.8000 202.0000 30.4000 ;
	    RECT 190.0000 26.8000 190.8000 28.4000 ;
	    RECT 195.4000 28.2000 197.0000 28.4000 ;
	    RECT 195.2000 27.8000 197.0000 28.2000 ;
	    RECT 180.4000 26.0000 184.4000 26.2000 ;
	    RECT 180.4000 22.2000 181.2000 26.0000 ;
	    RECT 183.6000 22.2000 184.4000 26.0000 ;
	    RECT 185.2000 22.2000 186.0000 26.2000 ;
	    RECT 187.4000 25.6000 189.2000 26.2000 ;
	    RECT 187.4000 24.4000 188.2000 25.6000 ;
	    RECT 187.4000 23.6000 189.2000 24.4000 ;
	    RECT 187.4000 22.2000 188.2000 23.6000 ;
	    RECT 195.2000 22.2000 196.0000 27.8000 ;
	    RECT 198.0000 27.6000 200.6000 28.4000 ;
	    RECT 198.2000 26.2000 198.8000 27.6000 ;
	    RECT 199.8000 26.2000 203.4000 26.6000 ;
	    RECT 198.0000 22.2000 198.8000 26.2000 ;
	    RECT 199.6000 26.0000 203.6000 26.2000 ;
	    RECT 199.6000 22.2000 200.4000 26.0000 ;
	    RECT 202.8000 22.2000 203.6000 26.0000 ;
	    RECT 204.4000 24.8000 205.2000 26.4000 ;
	    RECT 206.0000 22.2000 206.8000 31.7000 ;
	    RECT 207.6000 31.6000 208.4000 31.7000 ;
	    RECT 209.6000 28.4000 210.2000 31.8000 ;
	    RECT 210.8000 28.8000 211.6000 30.4000 ;
	    RECT 214.0000 30.3000 214.8000 32.4000 ;
	    RECT 212.5000 29.7000 214.8000 30.3000 ;
	    RECT 218.8000 31.6000 219.6000 32.4000 ;
	    RECT 222.0000 31.8000 223.8000 32.6000 ;
	    RECT 212.5000 28.4000 213.1000 29.7000 ;
	    RECT 218.8000 28.4000 219.4000 31.6000 ;
	    RECT 222.2000 28.4000 222.8000 31.8000 ;
	    RECT 207.6000 27.6000 210.2000 28.4000 ;
	    RECT 212.4000 28.2000 213.2000 28.4000 ;
	    RECT 217.8000 28.2000 219.4000 28.4000 ;
	    RECT 211.6000 27.6000 213.2000 28.2000 ;
	    RECT 217.6000 27.8000 219.4000 28.2000 ;
	    RECT 207.8000 26.2000 208.4000 27.6000 ;
	    RECT 211.6000 27.2000 212.4000 27.6000 ;
	    RECT 209.4000 26.2000 213.0000 26.6000 ;
	    RECT 207.6000 22.2000 208.4000 26.2000 ;
	    RECT 209.2000 26.0000 213.2000 26.2000 ;
	    RECT 209.2000 22.2000 210.0000 26.0000 ;
	    RECT 212.4000 22.2000 213.2000 26.0000 ;
	    RECT 217.6000 22.2000 218.4000 27.8000 ;
	    RECT 222.0000 27.6000 222.8000 28.4000 ;
	    RECT 222.2000 24.2000 222.8000 27.6000 ;
	    RECT 222.0000 22.2000 222.8000 24.2000 ;
	    RECT 4.4000 15.2000 5.2000 19.8000 ;
	    RECT 7.6000 16.0000 8.4000 19.8000 ;
	    RECT 3.0000 14.6000 5.2000 15.2000 ;
	    RECT 7.4000 15.2000 8.4000 16.0000 ;
	    RECT 3.0000 11.6000 3.6000 14.6000 ;
	    RECT 4.4000 12.3000 5.2000 13.2000 ;
	    RECT 7.4000 12.3000 8.2000 15.2000 ;
	    RECT 9.2000 14.6000 10.0000 19.8000 ;
	    RECT 15.6000 16.6000 16.4000 19.8000 ;
	    RECT 17.2000 17.0000 18.0000 19.8000 ;
	    RECT 18.8000 17.0000 19.6000 19.8000 ;
	    RECT 20.4000 17.0000 21.2000 19.8000 ;
	    RECT 22.0000 17.0000 22.8000 19.8000 ;
	    RECT 25.2000 17.0000 26.0000 19.8000 ;
	    RECT 28.4000 17.0000 29.2000 19.8000 ;
	    RECT 30.0000 17.0000 30.8000 19.8000 ;
	    RECT 31.6000 17.0000 32.4000 19.8000 ;
	    RECT 14.0000 15.8000 16.4000 16.6000 ;
	    RECT 33.2000 16.6000 34.0000 19.8000 ;
	    RECT 14.0000 15.2000 14.8000 15.8000 ;
	    RECT 4.4000 11.7000 8.2000 12.3000 ;
	    RECT 4.4000 11.6000 5.2000 11.7000 ;
	    RECT 2.4000 10.8000 3.6000 11.6000 ;
	    RECT 3.0000 10.2000 3.6000 10.8000 ;
	    RECT 7.4000 10.8000 8.2000 11.7000 ;
	    RECT 8.8000 14.0000 10.0000 14.6000 ;
	    RECT 13.0000 14.6000 14.8000 15.2000 ;
	    RECT 18.8000 15.6000 19.8000 16.4000 ;
	    RECT 22.8000 15.6000 24.4000 16.4000 ;
	    RECT 25.2000 15.8000 29.8000 16.4000 ;
	    RECT 33.2000 15.8000 35.8000 16.6000 ;
	    RECT 25.2000 15.6000 26.0000 15.8000 ;
	    RECT 8.8000 12.0000 9.4000 14.0000 ;
	    RECT 13.0000 13.4000 13.8000 14.6000 ;
	    RECT 10.0000 12.6000 13.8000 13.4000 ;
	    RECT 18.8000 12.8000 19.6000 15.6000 ;
	    RECT 25.2000 14.8000 26.0000 15.0000 ;
	    RECT 21.6000 14.2000 26.0000 14.8000 ;
	    RECT 21.6000 14.0000 22.4000 14.2000 ;
	    RECT 26.8000 13.6000 27.6000 15.2000 ;
	    RECT 29.0000 13.4000 29.8000 15.8000 ;
	    RECT 35.0000 15.2000 35.8000 15.8000 ;
	    RECT 35.0000 14.4000 38.0000 15.2000 ;
	    RECT 39.6000 13.8000 40.4000 19.8000 ;
	    RECT 22.0000 12.6000 25.2000 13.4000 ;
	    RECT 29.0000 12.6000 31.0000 13.4000 ;
	    RECT 31.6000 13.0000 40.4000 13.8000 ;
	    RECT 15.6000 12.0000 16.4000 12.6000 ;
	    RECT 33.2000 12.0000 34.0000 12.4000 ;
	    RECT 34.8000 12.0000 35.6000 12.4000 ;
	    RECT 36.4000 12.0000 37.2000 12.4000 ;
	    RECT 38.2000 12.0000 39.0000 12.2000 ;
	    RECT 8.8000 11.4000 9.6000 12.0000 ;
	    RECT 15.6000 11.4000 39.0000 12.0000 ;
	    RECT 3.0000 9.6000 5.2000 10.2000 ;
	    RECT 7.4000 10.0000 8.4000 10.8000 ;
	    RECT 4.4000 2.2000 5.2000 9.6000 ;
	    RECT 7.6000 2.2000 8.4000 10.0000 ;
	    RECT 9.0000 9.6000 9.6000 11.4000 ;
	    RECT 9.0000 9.0000 18.0000 9.6000 ;
	    RECT 9.0000 7.4000 9.6000 9.0000 ;
	    RECT 17.2000 8.8000 18.0000 9.0000 ;
	    RECT 20.4000 9.0000 29.0000 9.6000 ;
	    RECT 20.4000 8.8000 21.2000 9.0000 ;
	    RECT 12.2000 7.6000 14.8000 8.4000 ;
	    RECT 9.0000 6.8000 11.6000 7.4000 ;
	    RECT 10.8000 2.2000 11.6000 6.8000 ;
	    RECT 14.0000 2.2000 14.8000 7.6000 ;
	    RECT 15.4000 6.8000 19.6000 7.6000 ;
	    RECT 17.2000 2.2000 18.0000 5.0000 ;
	    RECT 18.8000 2.2000 19.6000 5.0000 ;
	    RECT 20.4000 2.2000 21.2000 5.0000 ;
	    RECT 22.0000 2.2000 22.8000 8.4000 ;
	    RECT 25.2000 7.6000 27.8000 8.4000 ;
	    RECT 28.4000 8.2000 29.0000 9.0000 ;
	    RECT 30.0000 9.4000 30.8000 9.6000 ;
	    RECT 30.0000 9.0000 35.4000 9.4000 ;
	    RECT 30.0000 8.8000 36.2000 9.0000 ;
	    RECT 34.8000 8.2000 36.2000 8.8000 ;
	    RECT 28.4000 7.6000 34.2000 8.2000 ;
	    RECT 37.2000 8.0000 38.8000 8.8000 ;
	    RECT 37.2000 7.6000 37.8000 8.0000 ;
	    RECT 25.2000 2.2000 26.0000 7.0000 ;
	    RECT 28.4000 2.2000 29.2000 7.0000 ;
	    RECT 33.6000 6.8000 37.8000 7.6000 ;
	    RECT 39.6000 7.4000 40.4000 13.0000 ;
	    RECT 38.4000 6.8000 40.4000 7.4000 ;
	    RECT 41.2000 13.8000 42.0000 19.8000 ;
	    RECT 47.6000 16.6000 48.4000 19.8000 ;
	    RECT 49.2000 17.0000 50.0000 19.8000 ;
	    RECT 50.8000 17.0000 51.6000 19.8000 ;
	    RECT 52.4000 17.0000 53.2000 19.8000 ;
	    RECT 55.6000 17.0000 56.4000 19.8000 ;
	    RECT 58.8000 17.0000 59.6000 19.8000 ;
	    RECT 60.4000 17.0000 61.2000 19.8000 ;
	    RECT 62.0000 17.0000 62.8000 19.8000 ;
	    RECT 63.6000 17.0000 64.4000 19.8000 ;
	    RECT 45.8000 15.8000 48.4000 16.6000 ;
	    RECT 65.2000 16.6000 66.0000 19.8000 ;
	    RECT 51.8000 15.8000 56.4000 16.4000 ;
	    RECT 45.8000 15.2000 46.6000 15.8000 ;
	    RECT 43.6000 14.4000 46.6000 15.2000 ;
	    RECT 41.2000 13.0000 50.0000 13.8000 ;
	    RECT 51.8000 13.4000 52.6000 15.8000 ;
	    RECT 55.6000 15.6000 56.4000 15.8000 ;
	    RECT 57.2000 15.6000 58.8000 16.4000 ;
	    RECT 61.8000 15.6000 62.8000 16.4000 ;
	    RECT 65.2000 15.8000 67.6000 16.6000 ;
	    RECT 54.0000 13.6000 54.8000 15.2000 ;
	    RECT 55.6000 14.8000 56.4000 15.0000 ;
	    RECT 55.6000 14.2000 60.0000 14.8000 ;
	    RECT 59.2000 14.0000 60.0000 14.2000 ;
	    RECT 41.2000 7.4000 42.0000 13.0000 ;
	    RECT 50.6000 12.6000 52.6000 13.4000 ;
	    RECT 56.4000 12.6000 59.6000 13.4000 ;
	    RECT 62.0000 12.8000 62.8000 15.6000 ;
	    RECT 66.8000 15.2000 67.6000 15.8000 ;
	    RECT 66.8000 14.6000 68.6000 15.2000 ;
	    RECT 67.8000 13.4000 68.6000 14.6000 ;
	    RECT 71.6000 14.6000 72.4000 19.8000 ;
	    RECT 73.2000 16.0000 74.0000 19.8000 ;
	    RECT 73.2000 15.2000 74.2000 16.0000 ;
	    RECT 71.6000 14.0000 72.8000 14.6000 ;
	    RECT 67.8000 12.6000 71.6000 13.4000 ;
	    RECT 42.6000 12.0000 43.4000 12.2000 ;
	    RECT 44.4000 12.0000 45.2000 12.4000 ;
	    RECT 47.6000 12.0000 48.4000 12.4000 ;
	    RECT 65.2000 12.0000 66.0000 12.6000 ;
	    RECT 72.2000 12.0000 72.8000 14.0000 ;
	    RECT 42.6000 11.4000 66.0000 12.0000 ;
	    RECT 72.0000 11.4000 72.8000 12.0000 ;
	    RECT 73.4000 12.3000 74.2000 15.2000 ;
	    RECT 81.2000 15.2000 82.0000 19.8000 ;
	    RECT 89.2000 15.2000 90.0000 19.8000 ;
	    RECT 92.4000 16.0000 93.2000 19.8000 ;
	    RECT 81.2000 14.6000 83.4000 15.2000 ;
	    RECT 81.2000 12.3000 82.0000 13.2000 ;
	    RECT 73.4000 11.7000 82.0000 12.3000 ;
	    RECT 72.0000 9.6000 72.6000 11.4000 ;
	    RECT 73.4000 10.8000 74.2000 11.7000 ;
	    RECT 81.2000 11.6000 82.0000 11.7000 ;
	    RECT 82.8000 11.6000 83.4000 14.6000 ;
	    RECT 87.8000 14.6000 90.0000 15.2000 ;
	    RECT 92.2000 15.2000 93.2000 16.0000 ;
	    RECT 87.8000 11.6000 88.4000 14.6000 ;
	    RECT 89.2000 12.3000 90.0000 13.2000 ;
	    RECT 92.2000 12.3000 93.0000 15.2000 ;
	    RECT 94.0000 14.6000 94.8000 19.8000 ;
	    RECT 100.4000 16.6000 101.2000 19.8000 ;
	    RECT 102.0000 17.0000 102.8000 19.8000 ;
	    RECT 103.6000 17.0000 104.4000 19.8000 ;
	    RECT 105.2000 17.0000 106.0000 19.8000 ;
	    RECT 106.8000 17.0000 107.6000 19.8000 ;
	    RECT 110.0000 17.0000 110.8000 19.8000 ;
	    RECT 113.2000 17.0000 114.0000 19.8000 ;
	    RECT 114.8000 17.0000 115.6000 19.8000 ;
	    RECT 116.4000 17.0000 117.2000 19.8000 ;
	    RECT 98.8000 15.8000 101.2000 16.6000 ;
	    RECT 118.0000 16.6000 118.8000 19.8000 ;
	    RECT 98.8000 15.2000 99.6000 15.8000 ;
	    RECT 89.2000 11.7000 93.0000 12.3000 ;
	    RECT 89.2000 11.6000 90.0000 11.7000 ;
	    RECT 50.8000 9.4000 51.6000 9.6000 ;
	    RECT 46.2000 9.0000 51.6000 9.4000 ;
	    RECT 45.4000 8.8000 51.6000 9.0000 ;
	    RECT 52.6000 9.0000 61.2000 9.6000 ;
	    RECT 42.8000 8.0000 44.4000 8.8000 ;
	    RECT 45.4000 8.2000 46.8000 8.8000 ;
	    RECT 52.6000 8.2000 53.2000 9.0000 ;
	    RECT 60.4000 8.8000 61.2000 9.0000 ;
	    RECT 63.6000 9.0000 72.6000 9.6000 ;
	    RECT 63.6000 8.8000 64.4000 9.0000 ;
	    RECT 43.8000 7.6000 44.4000 8.0000 ;
	    RECT 47.4000 7.6000 53.2000 8.2000 ;
	    RECT 53.8000 7.6000 56.4000 8.4000 ;
	    RECT 41.2000 6.8000 43.2000 7.4000 ;
	    RECT 43.8000 6.8000 48.0000 7.6000 ;
	    RECT 30.0000 2.2000 30.8000 5.0000 ;
	    RECT 31.6000 2.2000 32.4000 5.0000 ;
	    RECT 34.8000 2.2000 35.6000 6.8000 ;
	    RECT 38.4000 6.2000 39.0000 6.8000 ;
	    RECT 38.0000 5.6000 39.0000 6.2000 ;
	    RECT 42.6000 6.2000 43.2000 6.8000 ;
	    RECT 42.6000 5.6000 43.6000 6.2000 ;
	    RECT 38.0000 2.2000 38.8000 5.6000 ;
	    RECT 42.8000 2.2000 43.6000 5.6000 ;
	    RECT 46.0000 2.2000 46.8000 6.8000 ;
	    RECT 49.2000 2.2000 50.0000 5.0000 ;
	    RECT 50.8000 2.2000 51.6000 5.0000 ;
	    RECT 52.4000 2.2000 53.2000 7.0000 ;
	    RECT 55.6000 2.2000 56.4000 7.0000 ;
	    RECT 58.8000 2.2000 59.6000 8.4000 ;
	    RECT 66.8000 7.6000 69.4000 8.4000 ;
	    RECT 62.0000 6.8000 66.2000 7.6000 ;
	    RECT 60.4000 2.2000 61.2000 5.0000 ;
	    RECT 62.0000 2.2000 62.8000 5.0000 ;
	    RECT 63.6000 2.2000 64.4000 5.0000 ;
	    RECT 66.8000 2.2000 67.6000 7.6000 ;
	    RECT 72.0000 7.4000 72.6000 9.0000 ;
	    RECT 70.0000 6.8000 72.6000 7.4000 ;
	    RECT 73.2000 10.0000 74.2000 10.8000 ;
	    RECT 82.8000 10.8000 84.0000 11.6000 ;
	    RECT 87.2000 10.8000 88.4000 11.6000 ;
	    RECT 82.8000 10.2000 83.4000 10.8000 ;
	    RECT 70.0000 2.2000 70.8000 6.8000 ;
	    RECT 73.2000 2.2000 74.0000 10.0000 ;
	    RECT 81.2000 9.6000 83.4000 10.2000 ;
	    RECT 87.8000 10.2000 88.4000 10.8000 ;
	    RECT 92.2000 10.8000 93.0000 11.7000 ;
	    RECT 93.6000 14.0000 94.8000 14.6000 ;
	    RECT 97.8000 14.6000 99.6000 15.2000 ;
	    RECT 103.6000 15.6000 104.6000 16.4000 ;
	    RECT 107.6000 15.6000 109.2000 16.4000 ;
	    RECT 110.0000 15.8000 114.6000 16.4000 ;
	    RECT 118.0000 15.8000 120.6000 16.6000 ;
	    RECT 110.0000 15.6000 110.8000 15.8000 ;
	    RECT 93.6000 12.0000 94.2000 14.0000 ;
	    RECT 97.8000 13.4000 98.6000 14.6000 ;
	    RECT 94.8000 12.6000 98.6000 13.4000 ;
	    RECT 103.6000 12.8000 104.4000 15.6000 ;
	    RECT 110.0000 14.8000 110.8000 15.0000 ;
	    RECT 106.4000 14.2000 110.8000 14.8000 ;
	    RECT 106.4000 14.0000 107.2000 14.2000 ;
	    RECT 111.6000 13.6000 112.4000 15.2000 ;
	    RECT 113.8000 13.4000 114.6000 15.8000 ;
	    RECT 119.8000 15.2000 120.6000 15.8000 ;
	    RECT 119.8000 14.4000 122.8000 15.2000 ;
	    RECT 124.4000 13.8000 125.2000 19.8000 ;
	    RECT 126.0000 15.2000 126.8000 19.8000 ;
	    RECT 130.8000 15.2000 131.6000 19.8000 ;
	    RECT 137.2000 17.6000 138.0000 19.8000 ;
	    RECT 135.6000 15.6000 136.4000 17.2000 ;
	    RECT 126.0000 14.6000 128.2000 15.2000 ;
	    RECT 130.8000 14.6000 133.0000 15.2000 ;
	    RECT 106.8000 12.6000 110.0000 13.4000 ;
	    RECT 113.8000 12.6000 115.8000 13.4000 ;
	    RECT 116.4000 13.0000 125.2000 13.8000 ;
	    RECT 100.4000 12.0000 101.2000 12.6000 ;
	    RECT 118.0000 12.0000 118.8000 12.4000 ;
	    RECT 121.2000 12.0000 122.0000 12.4000 ;
	    RECT 123.0000 12.0000 123.8000 12.2000 ;
	    RECT 93.6000 11.4000 94.4000 12.0000 ;
	    RECT 100.4000 11.4000 123.8000 12.0000 ;
	    RECT 87.8000 9.6000 90.0000 10.2000 ;
	    RECT 92.2000 10.0000 93.2000 10.8000 ;
	    RECT 81.2000 2.2000 82.0000 9.6000 ;
	    RECT 89.2000 2.2000 90.0000 9.6000 ;
	    RECT 92.4000 2.2000 93.2000 10.0000 ;
	    RECT 93.8000 9.6000 94.4000 11.4000 ;
	    RECT 93.8000 9.0000 102.8000 9.6000 ;
	    RECT 93.8000 7.4000 94.4000 9.0000 ;
	    RECT 102.0000 8.8000 102.8000 9.0000 ;
	    RECT 105.2000 9.0000 113.8000 9.6000 ;
	    RECT 105.2000 8.8000 106.0000 9.0000 ;
	    RECT 97.0000 7.6000 99.6000 8.4000 ;
	    RECT 93.8000 6.8000 96.4000 7.4000 ;
	    RECT 95.6000 2.2000 96.4000 6.8000 ;
	    RECT 98.8000 2.2000 99.6000 7.6000 ;
	    RECT 100.2000 6.8000 104.4000 7.6000 ;
	    RECT 102.0000 2.2000 102.8000 5.0000 ;
	    RECT 103.6000 2.2000 104.4000 5.0000 ;
	    RECT 105.2000 2.2000 106.0000 5.0000 ;
	    RECT 106.8000 2.2000 107.6000 8.4000 ;
	    RECT 110.0000 7.6000 112.6000 8.4000 ;
	    RECT 113.2000 8.2000 113.8000 9.0000 ;
	    RECT 114.8000 9.4000 115.6000 9.6000 ;
	    RECT 114.8000 9.0000 120.2000 9.4000 ;
	    RECT 114.8000 8.8000 121.0000 9.0000 ;
	    RECT 119.6000 8.2000 121.0000 8.8000 ;
	    RECT 113.2000 7.6000 119.0000 8.2000 ;
	    RECT 122.0000 8.0000 123.6000 8.8000 ;
	    RECT 122.0000 7.6000 122.6000 8.0000 ;
	    RECT 110.0000 2.2000 110.8000 7.0000 ;
	    RECT 113.2000 2.2000 114.0000 7.0000 ;
	    RECT 118.4000 6.8000 122.6000 7.6000 ;
	    RECT 124.4000 7.4000 125.2000 13.0000 ;
	    RECT 126.0000 11.6000 126.8000 13.2000 ;
	    RECT 127.6000 11.6000 128.2000 14.6000 ;
	    RECT 130.8000 11.6000 131.6000 13.2000 ;
	    RECT 132.4000 11.6000 133.0000 14.6000 ;
	    RECT 137.4000 14.4000 138.0000 17.6000 ;
	    RECT 140.4000 15.8000 141.2000 19.8000 ;
	    RECT 144.6000 16.8000 145.4000 19.8000 ;
	    RECT 144.6000 15.8000 146.0000 16.8000 ;
	    RECT 146.8000 16.0000 147.6000 19.8000 ;
	    RECT 150.0000 16.0000 150.8000 19.8000 ;
	    RECT 146.8000 15.8000 150.8000 16.0000 ;
	    RECT 151.6000 15.8000 152.4000 19.8000 ;
	    RECT 140.6000 15.6000 141.2000 15.8000 ;
	    RECT 140.6000 15.2000 142.4000 15.6000 ;
	    RECT 140.6000 15.0000 144.8000 15.2000 ;
	    RECT 141.8000 14.6000 144.8000 15.0000 ;
	    RECT 144.0000 14.4000 144.8000 14.6000 ;
	    RECT 137.2000 13.6000 138.0000 14.4000 ;
	    RECT 127.6000 10.8000 128.8000 11.6000 ;
	    RECT 132.4000 10.8000 133.6000 11.6000 ;
	    RECT 127.6000 10.2000 128.2000 10.8000 ;
	    RECT 132.4000 10.2000 133.0000 10.8000 ;
	    RECT 137.4000 10.2000 138.0000 13.6000 ;
	    RECT 138.8000 12.3000 139.6000 12.4000 ;
	    RECT 140.4000 12.3000 141.2000 14.4000 ;
	    RECT 142.4000 13.8000 143.2000 14.0000 ;
	    RECT 142.2000 13.2000 143.2000 13.8000 ;
	    RECT 142.2000 12.4000 142.8000 13.2000 ;
	    RECT 138.8000 11.7000 141.2000 12.3000 ;
	    RECT 138.8000 10.8000 139.6000 11.7000 ;
	    RECT 142.0000 11.6000 142.8000 12.4000 ;
	    RECT 144.0000 11.0000 144.6000 14.4000 ;
	    RECT 145.4000 12.4000 146.0000 15.8000 ;
	    RECT 147.0000 15.4000 150.6000 15.8000 ;
	    RECT 147.6000 14.4000 148.4000 14.8000 ;
	    RECT 151.6000 14.4000 152.2000 15.8000 ;
	    RECT 153.2000 15.6000 154.0000 19.8000 ;
	    RECT 154.8000 16.0000 155.6000 19.8000 ;
	    RECT 158.0000 16.0000 158.8000 19.8000 ;
	    RECT 154.8000 15.8000 158.8000 16.0000 ;
	    RECT 153.4000 14.4000 154.0000 15.6000 ;
	    RECT 155.0000 15.4000 158.6000 15.8000 ;
	    RECT 167.6000 15.2000 168.4000 19.8000 ;
	    RECT 169.2000 16.3000 170.0000 16.4000 ;
	    RECT 170.8000 16.3000 171.6000 19.8000 ;
	    RECT 169.2000 15.7000 171.6000 16.3000 ;
	    RECT 169.2000 15.6000 170.0000 15.7000 ;
	    RECT 157.2000 14.4000 158.0000 14.8000 ;
	    RECT 166.2000 14.6000 168.4000 15.2000 ;
	    RECT 170.6000 15.2000 171.6000 15.7000 ;
	    RECT 146.8000 13.8000 148.4000 14.4000 ;
	    RECT 146.8000 13.6000 147.6000 13.8000 ;
	    RECT 149.8000 13.6000 152.4000 14.4000 ;
	    RECT 153.2000 13.6000 155.8000 14.4000 ;
	    RECT 157.2000 14.3000 158.8000 14.4000 ;
	    RECT 161.2000 14.3000 162.0000 14.4000 ;
	    RECT 157.2000 13.8000 162.0000 14.3000 ;
	    RECT 158.0000 13.7000 162.0000 13.8000 ;
	    RECT 158.0000 13.6000 158.8000 13.7000 ;
	    RECT 161.2000 13.6000 162.0000 13.7000 ;
	    RECT 145.2000 12.3000 146.0000 12.4000 ;
	    RECT 148.4000 12.3000 149.2000 13.2000 ;
	    RECT 145.2000 11.7000 149.2000 12.3000 ;
	    RECT 145.2000 11.6000 146.0000 11.7000 ;
	    RECT 148.4000 11.6000 149.2000 11.7000 ;
	    RECT 149.8000 12.3000 150.4000 13.6000 ;
	    RECT 149.8000 11.7000 153.9000 12.3000 ;
	    RECT 142.2000 10.4000 144.6000 11.0000 ;
	    RECT 123.2000 6.8000 125.2000 7.4000 ;
	    RECT 126.0000 9.6000 128.2000 10.2000 ;
	    RECT 130.8000 9.6000 133.0000 10.2000 ;
	    RECT 114.8000 2.2000 115.6000 5.0000 ;
	    RECT 116.4000 2.2000 117.2000 5.0000 ;
	    RECT 119.6000 2.2000 120.4000 6.8000 ;
	    RECT 123.2000 6.2000 123.8000 6.8000 ;
	    RECT 122.8000 5.6000 123.8000 6.2000 ;
	    RECT 122.8000 2.2000 123.6000 5.6000 ;
	    RECT 126.0000 2.2000 126.8000 9.6000 ;
	    RECT 130.8000 2.2000 131.6000 9.6000 ;
	    RECT 137.2000 9.4000 139.0000 10.2000 ;
	    RECT 138.2000 2.2000 139.0000 9.4000 ;
	    RECT 142.2000 6.2000 142.8000 10.4000 ;
	    RECT 145.4000 10.2000 146.0000 11.6000 ;
	    RECT 149.8000 10.2000 150.4000 11.7000 ;
	    RECT 153.3000 10.4000 153.9000 11.7000 ;
	    RECT 151.6000 10.2000 152.4000 10.4000 ;
	    RECT 142.0000 2.2000 142.8000 6.2000 ;
	    RECT 145.2000 2.2000 146.0000 10.2000 ;
	    RECT 149.4000 9.6000 150.4000 10.2000 ;
	    RECT 151.0000 9.6000 152.4000 10.2000 ;
	    RECT 153.2000 10.2000 154.0000 10.4000 ;
	    RECT 155.2000 10.2000 155.8000 13.6000 ;
	    RECT 156.4000 11.6000 157.2000 13.2000 ;
	    RECT 166.2000 11.6000 166.8000 14.6000 ;
	    RECT 167.6000 12.3000 168.4000 13.2000 ;
	    RECT 170.6000 12.3000 171.4000 15.2000 ;
	    RECT 172.4000 14.6000 173.2000 19.8000 ;
	    RECT 178.8000 16.6000 179.6000 19.8000 ;
	    RECT 180.4000 17.0000 181.2000 19.8000 ;
	    RECT 182.0000 17.0000 182.8000 19.8000 ;
	    RECT 183.6000 17.0000 184.4000 19.8000 ;
	    RECT 185.2000 17.0000 186.0000 19.8000 ;
	    RECT 188.4000 17.0000 189.2000 19.8000 ;
	    RECT 191.6000 17.0000 192.4000 19.8000 ;
	    RECT 193.2000 17.0000 194.0000 19.8000 ;
	    RECT 194.8000 17.0000 195.6000 19.8000 ;
	    RECT 177.2000 15.8000 179.6000 16.6000 ;
	    RECT 196.4000 16.6000 197.2000 19.8000 ;
	    RECT 177.2000 15.2000 178.0000 15.8000 ;
	    RECT 167.6000 11.7000 171.4000 12.3000 ;
	    RECT 167.6000 11.6000 168.4000 11.7000 ;
	    RECT 165.6000 10.8000 166.8000 11.6000 ;
	    RECT 166.2000 10.2000 166.8000 10.8000 ;
	    RECT 170.6000 10.8000 171.4000 11.7000 ;
	    RECT 172.0000 14.0000 173.2000 14.6000 ;
	    RECT 176.2000 14.6000 178.0000 15.2000 ;
	    RECT 182.0000 15.6000 183.0000 16.4000 ;
	    RECT 186.0000 15.6000 187.6000 16.4000 ;
	    RECT 188.4000 15.8000 193.0000 16.4000 ;
	    RECT 196.4000 15.8000 199.0000 16.6000 ;
	    RECT 188.4000 15.6000 189.2000 15.8000 ;
	    RECT 172.0000 12.0000 172.6000 14.0000 ;
	    RECT 176.2000 13.4000 177.0000 14.6000 ;
	    RECT 173.2000 12.6000 177.0000 13.4000 ;
	    RECT 182.0000 12.8000 182.8000 15.6000 ;
	    RECT 188.4000 14.8000 189.2000 15.0000 ;
	    RECT 184.8000 14.2000 189.2000 14.8000 ;
	    RECT 184.8000 14.0000 185.6000 14.2000 ;
	    RECT 190.0000 13.6000 190.8000 15.2000 ;
	    RECT 192.2000 13.4000 193.0000 15.8000 ;
	    RECT 198.2000 15.2000 199.0000 15.8000 ;
	    RECT 198.2000 14.4000 201.2000 15.2000 ;
	    RECT 202.8000 13.8000 203.6000 19.8000 ;
	    RECT 204.4000 16.0000 205.2000 19.8000 ;
	    RECT 207.6000 16.0000 208.4000 19.8000 ;
	    RECT 204.4000 15.8000 208.4000 16.0000 ;
	    RECT 209.2000 15.8000 210.0000 19.8000 ;
	    RECT 204.6000 15.4000 208.2000 15.8000 ;
	    RECT 209.2000 14.4000 209.8000 15.8000 ;
	    RECT 185.2000 12.6000 188.4000 13.4000 ;
	    RECT 192.2000 12.6000 194.2000 13.4000 ;
	    RECT 194.8000 13.0000 203.6000 13.8000 ;
	    RECT 207.4000 13.6000 210.0000 14.4000 ;
	    RECT 178.8000 12.0000 179.6000 12.6000 ;
	    RECT 196.4000 12.0000 197.2000 12.4000 ;
	    RECT 201.4000 12.0000 202.2000 12.2000 ;
	    RECT 172.0000 11.4000 172.8000 12.0000 ;
	    RECT 178.8000 11.4000 202.2000 12.0000 ;
	    RECT 153.2000 9.6000 154.6000 10.2000 ;
	    RECT 155.2000 9.6000 156.2000 10.2000 ;
	    RECT 166.2000 9.6000 168.4000 10.2000 ;
	    RECT 170.6000 10.0000 171.6000 10.8000 ;
	    RECT 149.4000 2.2000 150.2000 9.6000 ;
	    RECT 151.0000 8.4000 151.6000 9.6000 ;
	    RECT 150.8000 7.6000 151.6000 8.4000 ;
	    RECT 154.0000 8.4000 154.6000 9.6000 ;
	    RECT 154.0000 7.6000 154.8000 8.4000 ;
	    RECT 155.4000 2.2000 156.2000 9.6000 ;
	    RECT 167.6000 2.2000 168.4000 9.6000 ;
	    RECT 170.8000 2.2000 171.6000 10.0000 ;
	    RECT 172.2000 9.6000 172.8000 11.4000 ;
	    RECT 172.2000 9.0000 181.2000 9.6000 ;
	    RECT 172.2000 7.4000 172.8000 9.0000 ;
	    RECT 180.4000 8.8000 181.2000 9.0000 ;
	    RECT 183.6000 9.0000 192.2000 9.6000 ;
	    RECT 183.6000 8.8000 184.4000 9.0000 ;
	    RECT 175.4000 7.6000 178.0000 8.4000 ;
	    RECT 172.2000 6.8000 174.8000 7.4000 ;
	    RECT 174.0000 2.2000 174.8000 6.8000 ;
	    RECT 177.2000 2.2000 178.0000 7.6000 ;
	    RECT 178.6000 6.8000 182.8000 7.6000 ;
	    RECT 180.4000 2.2000 181.2000 5.0000 ;
	    RECT 182.0000 2.2000 182.8000 5.0000 ;
	    RECT 183.6000 2.2000 184.4000 5.0000 ;
	    RECT 185.2000 2.2000 186.0000 8.4000 ;
	    RECT 188.4000 7.6000 191.0000 8.4000 ;
	    RECT 191.6000 8.2000 192.2000 9.0000 ;
	    RECT 193.2000 9.4000 194.0000 9.6000 ;
	    RECT 193.2000 9.0000 198.6000 9.4000 ;
	    RECT 193.2000 8.8000 199.4000 9.0000 ;
	    RECT 198.0000 8.2000 199.4000 8.8000 ;
	    RECT 191.6000 7.6000 197.4000 8.2000 ;
	    RECT 200.4000 8.0000 202.0000 8.8000 ;
	    RECT 200.4000 7.6000 201.0000 8.0000 ;
	    RECT 188.4000 2.2000 189.2000 7.0000 ;
	    RECT 191.6000 2.2000 192.4000 7.0000 ;
	    RECT 196.8000 6.8000 201.0000 7.6000 ;
	    RECT 202.8000 7.4000 203.6000 13.0000 ;
	    RECT 206.0000 11.6000 206.8000 13.2000 ;
	    RECT 207.4000 10.2000 208.0000 13.6000 ;
	    RECT 209.2000 10.2000 210.0000 10.4000 ;
	    RECT 201.6000 6.8000 203.6000 7.4000 ;
	    RECT 207.0000 9.6000 208.0000 10.2000 ;
	    RECT 208.6000 9.6000 210.0000 10.2000 ;
	    RECT 193.2000 2.2000 194.0000 5.0000 ;
	    RECT 194.8000 2.2000 195.6000 5.0000 ;
	    RECT 198.0000 2.2000 198.8000 6.8000 ;
	    RECT 201.6000 6.2000 202.2000 6.8000 ;
	    RECT 201.2000 5.6000 202.2000 6.2000 ;
	    RECT 201.2000 2.2000 202.0000 5.6000 ;
	    RECT 207.0000 2.2000 207.8000 9.6000 ;
	    RECT 208.6000 8.4000 209.2000 9.6000 ;
	    RECT 208.4000 7.6000 209.2000 8.4000 ;
	    RECT 210.8000 2.2000 211.6000 19.8000 ;
	    RECT 212.4000 10.3000 213.2000 10.4000 ;
	    RECT 214.0000 10.3000 214.8000 19.8000 ;
	    RECT 212.4000 9.7000 214.8000 10.3000 ;
	    RECT 212.4000 9.6000 213.2000 9.7000 ;
	    RECT 214.0000 2.2000 214.8000 9.7000 ;
	    RECT 217.2000 2.2000 218.0000 19.8000 ;
	    RECT 218.8000 15.6000 219.6000 17.2000 ;
	    RECT 220.4000 15.2000 221.2000 19.8000 ;
	    RECT 220.4000 14.6000 222.6000 15.2000 ;
	    RECT 220.4000 11.6000 221.2000 13.2000 ;
	    RECT 222.0000 11.6000 222.6000 14.6000 ;
	    RECT 222.0000 10.8000 223.2000 11.6000 ;
	    RECT 222.0000 10.2000 222.6000 10.8000 ;
	    RECT 220.4000 9.6000 222.6000 10.2000 ;
	    RECT 220.4000 2.2000 221.2000 9.6000 ;
         LAYER metal2 ;
	    RECT 14.0000 187.6000 14.8000 188.4000 ;
	    RECT 6.0000 185.6000 6.8000 186.4000 ;
	    RECT 6.1000 176.4000 6.7000 185.6000 ;
	    RECT 14.1000 178.4000 14.7000 187.6000 ;
	    RECT 17.2000 184.2000 18.0000 197.8000 ;
	    RECT 18.8000 184.2000 19.6000 197.8000 ;
	    RECT 20.4000 184.2000 21.2000 197.8000 ;
	    RECT 22.0000 184.2000 22.8000 195.8000 ;
	    RECT 23.6000 185.6000 24.4000 186.4000 ;
	    RECT 17.2000 181.6000 18.0000 182.4000 ;
	    RECT 14.0000 177.6000 14.8000 178.4000 ;
	    RECT 6.0000 175.6000 6.8000 176.4000 ;
	    RECT 17.3000 172.4000 17.9000 181.6000 ;
	    RECT 23.7000 176.4000 24.3000 185.6000 ;
	    RECT 25.2000 184.2000 26.0000 195.8000 ;
	    RECT 26.8000 187.6000 27.6000 188.4000 ;
	    RECT 28.4000 184.2000 29.2000 195.8000 ;
	    RECT 30.0000 184.2000 30.8000 197.8000 ;
	    RECT 31.6000 184.2000 32.4000 197.8000 ;
	    RECT 36.4000 189.6000 37.2000 190.4000 ;
	    RECT 36.5000 180.4000 37.1000 189.6000 ;
	    RECT 52.4000 183.6000 53.2000 184.4000 ;
	    RECT 57.2000 183.6000 58.0000 184.4000 ;
	    RECT 62.0000 184.2000 62.8000 197.8000 ;
	    RECT 63.6000 184.2000 64.4000 197.8000 ;
	    RECT 65.2000 184.2000 66.0000 197.8000 ;
	    RECT 66.8000 184.2000 67.6000 195.8000 ;
	    RECT 68.4000 185.6000 69.2000 186.4000 ;
	    RECT 36.4000 179.6000 37.2000 180.4000 ;
	    RECT 49.2000 179.6000 50.0000 180.4000 ;
	    RECT 23.6000 175.6000 24.4000 176.4000 ;
	    RECT 4.4000 171.6000 5.2000 172.4000 ;
	    RECT 15.6000 171.6000 16.4000 172.4000 ;
	    RECT 17.2000 171.6000 18.0000 172.4000 ;
	    RECT 4.5000 166.4000 5.1000 171.6000 ;
	    RECT 4.4000 165.6000 5.2000 166.4000 ;
	    RECT 14.0000 147.6000 14.8000 148.4000 ;
	    RECT 6.0000 145.6000 6.8000 146.4000 ;
	    RECT 4.4000 137.6000 5.2000 138.4000 ;
	    RECT 4.5000 132.4000 5.1000 137.6000 ;
	    RECT 6.1000 136.4000 6.7000 145.6000 ;
	    RECT 14.1000 138.4000 14.7000 147.6000 ;
	    RECT 14.0000 137.6000 14.8000 138.4000 ;
	    RECT 6.0000 135.6000 6.8000 136.4000 ;
	    RECT 15.7000 134.3000 16.3000 171.6000 ;
	    RECT 17.3000 160.4000 17.9000 171.6000 ;
	    RECT 20.4000 165.6000 21.2000 166.4000 ;
	    RECT 17.2000 159.6000 18.0000 160.4000 ;
	    RECT 17.2000 144.2000 18.0000 157.8000 ;
	    RECT 18.8000 144.2000 19.6000 157.8000 ;
	    RECT 20.4000 144.2000 21.2000 157.8000 ;
	    RECT 22.0000 144.2000 22.8000 155.8000 ;
	    RECT 23.7000 146.4000 24.3000 175.6000 ;
	    RECT 30.0000 164.2000 30.8000 177.8000 ;
	    RECT 31.6000 164.2000 32.4000 177.8000 ;
	    RECT 33.2000 164.2000 34.0000 177.8000 ;
	    RECT 34.8000 166.2000 35.6000 177.8000 ;
	    RECT 36.4000 175.6000 37.2000 176.4000 ;
	    RECT 38.0000 166.2000 38.8000 177.8000 ;
	    RECT 39.6000 177.6000 40.4000 178.4000 ;
	    RECT 39.7000 174.4000 40.3000 177.6000 ;
	    RECT 39.6000 173.6000 40.4000 174.4000 ;
	    RECT 39.6000 171.6000 40.4000 172.4000 ;
	    RECT 23.6000 145.6000 24.4000 146.4000 ;
	    RECT 25.2000 144.2000 26.0000 155.8000 ;
	    RECT 26.8000 147.6000 27.6000 148.4000 ;
	    RECT 28.4000 144.2000 29.2000 155.8000 ;
	    RECT 30.0000 144.2000 30.8000 157.8000 ;
	    RECT 31.6000 144.2000 32.4000 157.8000 ;
	    RECT 39.7000 150.4000 40.3000 171.6000 ;
	    RECT 41.2000 166.2000 42.0000 177.8000 ;
	    RECT 42.8000 164.2000 43.6000 177.8000 ;
	    RECT 44.4000 164.2000 45.2000 177.8000 ;
	    RECT 49.3000 172.4000 49.9000 179.6000 ;
	    RECT 57.3000 176.4000 57.9000 183.6000 ;
	    RECT 68.5000 176.4000 69.1000 185.6000 ;
	    RECT 70.0000 184.2000 70.8000 195.8000 ;
	    RECT 71.6000 187.6000 72.4000 188.4000 ;
	    RECT 71.7000 182.3000 72.3000 187.6000 ;
	    RECT 73.2000 184.2000 74.0000 195.8000 ;
	    RECT 74.8000 184.2000 75.6000 197.8000 ;
	    RECT 76.4000 184.2000 77.2000 197.8000 ;
	    RECT 81.2000 189.6000 82.0000 190.4000 ;
	    RECT 89.2000 189.6000 90.0000 190.4000 ;
	    RECT 90.8000 189.6000 91.6000 190.4000 ;
	    RECT 95.6000 189.6000 96.4000 190.4000 ;
	    RECT 100.4000 189.6000 101.2000 190.4000 ;
	    RECT 110.0000 189.6000 110.8000 190.4000 ;
	    RECT 118.0000 189.6000 118.8000 190.4000 ;
	    RECT 70.1000 181.7000 72.3000 182.3000 ;
	    RECT 70.1000 178.4000 70.7000 181.7000 ;
	    RECT 73.2000 181.6000 74.0000 182.4000 ;
	    RECT 70.0000 177.6000 70.8000 178.4000 ;
	    RECT 54.0000 175.6000 54.8000 176.4000 ;
	    RECT 57.2000 175.6000 58.0000 176.4000 ;
	    RECT 68.4000 175.6000 69.2000 176.4000 ;
	    RECT 49.2000 171.6000 50.0000 172.4000 ;
	    RECT 54.1000 166.4000 54.7000 175.6000 ;
	    RECT 73.3000 172.4000 73.9000 181.6000 ;
	    RECT 81.3000 180.4000 81.9000 189.6000 ;
	    RECT 81.2000 179.6000 82.0000 180.4000 ;
	    RECT 89.3000 178.4000 89.9000 189.6000 ;
	    RECT 90.9000 188.4000 91.5000 189.6000 ;
	    RECT 90.8000 187.6000 91.6000 188.4000 ;
	    RECT 78.0000 177.6000 78.8000 178.4000 ;
	    RECT 89.2000 177.6000 90.0000 178.4000 ;
	    RECT 79.6000 175.6000 80.4000 176.4000 ;
	    RECT 84.4000 175.6000 85.2000 176.4000 ;
	    RECT 84.5000 174.4000 85.1000 175.6000 ;
	    RECT 90.9000 174.4000 91.5000 187.6000 ;
	    RECT 76.4000 173.6000 77.2000 174.4000 ;
	    RECT 81.2000 173.6000 82.0000 174.4000 ;
	    RECT 84.4000 173.6000 85.2000 174.4000 ;
	    RECT 90.8000 173.6000 91.6000 174.4000 ;
	    RECT 57.2000 171.6000 58.0000 172.4000 ;
	    RECT 71.6000 171.6000 72.4000 172.4000 ;
	    RECT 73.2000 171.6000 74.0000 172.4000 ;
	    RECT 74.8000 171.6000 75.6000 172.4000 ;
	    RECT 82.8000 171.6000 83.6000 172.4000 ;
	    RECT 60.4000 167.6000 61.2000 168.4000 ;
	    RECT 54.0000 165.6000 54.8000 166.4000 ;
	    RECT 41.2000 151.6000 42.0000 152.4000 ;
	    RECT 36.4000 149.6000 37.2000 150.4000 ;
	    RECT 39.6000 149.6000 40.4000 150.4000 ;
	    RECT 41.3000 148.4000 41.9000 151.6000 ;
	    RECT 44.4000 149.6000 45.2000 150.4000 ;
	    RECT 52.4000 149.6000 53.2000 150.4000 ;
	    RECT 41.2000 147.6000 42.0000 148.4000 ;
	    RECT 42.8000 147.6000 43.6000 148.4000 ;
	    RECT 46.0000 147.6000 46.8000 148.4000 ;
	    RECT 42.9000 146.4000 43.5000 147.6000 ;
	    RECT 36.4000 145.6000 37.2000 146.4000 ;
	    RECT 42.8000 145.6000 43.6000 146.4000 ;
	    RECT 47.6000 145.6000 48.4000 146.4000 ;
	    RECT 20.4000 137.6000 21.2000 138.4000 ;
	    RECT 14.1000 133.7000 16.3000 134.3000 ;
	    RECT 4.4000 131.6000 5.2000 132.4000 ;
	    RECT 12.4000 121.6000 13.2000 122.4000 ;
	    RECT 12.5000 118.4000 13.1000 121.6000 ;
	    RECT 12.4000 117.6000 13.2000 118.4000 ;
	    RECT 14.1000 114.4000 14.7000 133.7000 ;
	    RECT 15.6000 131.6000 16.4000 132.4000 ;
	    RECT 17.2000 131.6000 18.0000 132.4000 ;
	    RECT 15.7000 122.4000 16.3000 131.6000 ;
	    RECT 28.4000 127.6000 29.2000 128.4000 ;
	    RECT 15.6000 121.6000 16.4000 122.4000 ;
	    RECT 14.0000 113.6000 14.8000 114.4000 ;
	    RECT 28.5000 112.4000 29.1000 127.6000 ;
	    RECT 30.0000 124.2000 30.8000 137.8000 ;
	    RECT 31.6000 124.2000 32.4000 137.8000 ;
	    RECT 33.2000 124.2000 34.0000 137.8000 ;
	    RECT 34.8000 126.2000 35.6000 137.8000 ;
	    RECT 36.5000 136.4000 37.1000 145.6000 ;
	    RECT 49.2000 143.6000 50.0000 144.4000 ;
	    RECT 36.4000 135.6000 37.2000 136.4000 ;
	    RECT 36.5000 124.4000 37.1000 135.6000 ;
	    RECT 38.0000 126.2000 38.8000 137.8000 ;
	    RECT 39.6000 133.6000 40.4000 134.4000 ;
	    RECT 41.2000 126.2000 42.0000 137.8000 ;
	    RECT 36.4000 123.6000 37.2000 124.4000 ;
	    RECT 42.8000 124.2000 43.6000 137.8000 ;
	    RECT 44.4000 124.2000 45.2000 137.8000 ;
	    RECT 49.3000 134.4000 49.9000 143.6000 ;
	    RECT 49.2000 133.6000 50.0000 134.4000 ;
	    RECT 52.5000 132.4000 53.1000 149.6000 ;
	    RECT 54.1000 148.4000 54.7000 165.6000 ;
	    RECT 60.5000 158.4000 61.1000 167.6000 ;
	    RECT 60.4000 157.6000 61.2000 158.4000 ;
	    RECT 54.0000 147.6000 54.8000 148.4000 ;
	    RECT 54.0000 145.6000 54.8000 146.4000 ;
	    RECT 54.1000 138.4000 54.7000 145.6000 ;
	    RECT 70.0000 144.2000 70.8000 157.8000 ;
	    RECT 71.6000 144.2000 72.4000 157.8000 ;
	    RECT 73.2000 144.2000 74.0000 155.8000 ;
	    RECT 74.9000 150.4000 75.5000 171.6000 ;
	    RECT 87.6000 169.6000 88.4000 170.4000 ;
	    RECT 74.8000 149.6000 75.6000 150.4000 ;
	    RECT 74.8000 147.6000 75.6000 148.4000 ;
	    RECT 74.9000 142.4000 75.5000 147.6000 ;
	    RECT 76.4000 144.2000 77.2000 155.8000 ;
	    RECT 78.0000 145.6000 78.8000 146.4000 ;
	    RECT 74.8000 141.6000 75.6000 142.4000 ;
	    RECT 78.1000 142.3000 78.7000 145.6000 ;
	    RECT 79.6000 144.2000 80.4000 155.8000 ;
	    RECT 81.2000 144.2000 82.0000 157.8000 ;
	    RECT 82.8000 144.2000 83.6000 157.8000 ;
	    RECT 84.4000 144.2000 85.2000 157.8000 ;
	    RECT 86.0000 149.6000 86.8000 150.4000 ;
	    RECT 76.5000 141.7000 78.7000 142.3000 ;
	    RECT 54.0000 137.6000 54.8000 138.4000 ;
	    RECT 54.1000 134.4000 54.7000 137.6000 ;
	    RECT 58.8000 135.6000 59.6000 136.4000 ;
	    RECT 74.8000 135.6000 75.6000 136.4000 ;
	    RECT 54.0000 133.6000 54.8000 134.4000 ;
	    RECT 60.4000 133.6000 61.2000 134.4000 ;
	    RECT 74.8000 133.6000 75.6000 134.4000 ;
	    RECT 60.5000 132.4000 61.1000 133.6000 ;
	    RECT 46.0000 131.6000 46.8000 132.4000 ;
	    RECT 52.4000 131.6000 53.2000 132.4000 ;
	    RECT 55.6000 131.6000 56.4000 132.4000 ;
	    RECT 60.4000 131.6000 61.2000 132.4000 ;
	    RECT 70.0000 131.6000 70.8000 132.4000 ;
	    RECT 31.6000 121.6000 32.4000 122.4000 ;
	    RECT 17.2000 111.6000 18.0000 112.4000 ;
	    RECT 25.2000 111.6000 26.0000 112.4000 ;
	    RECT 28.4000 111.6000 29.2000 112.4000 ;
	    RECT 17.3000 110.4000 17.9000 111.6000 ;
	    RECT 25.3000 110.4000 25.9000 111.6000 ;
	    RECT 4.4000 109.6000 5.2000 110.4000 ;
	    RECT 10.8000 109.6000 11.6000 110.4000 ;
	    RECT 17.2000 109.6000 18.0000 110.4000 ;
	    RECT 25.2000 109.6000 26.0000 110.4000 ;
	    RECT 4.5000 106.4000 5.1000 109.6000 ;
	    RECT 10.9000 108.4000 11.5000 109.6000 ;
	    RECT 10.8000 107.6000 11.6000 108.4000 ;
	    RECT 22.0000 107.6000 22.8000 108.4000 ;
	    RECT 26.8000 107.6000 27.6000 108.4000 ;
	    RECT 10.9000 106.4000 11.5000 107.6000 ;
	    RECT 26.9000 106.4000 27.5000 107.6000 ;
	    RECT 4.4000 106.3000 5.2000 106.4000 ;
	    RECT 2.9000 105.7000 5.2000 106.3000 ;
	    RECT 2.9000 98.4000 3.5000 105.7000 ;
	    RECT 4.4000 105.6000 5.2000 105.7000 ;
	    RECT 10.8000 105.6000 11.6000 106.4000 ;
	    RECT 14.0000 105.6000 14.8000 106.4000 ;
	    RECT 22.0000 105.6000 22.8000 106.4000 ;
	    RECT 26.8000 105.6000 27.6000 106.4000 ;
	    RECT 20.4000 103.6000 21.2000 104.4000 ;
	    RECT 20.5000 100.3000 21.1000 103.6000 ;
	    RECT 20.5000 99.7000 22.7000 100.3000 ;
	    RECT 2.8000 97.6000 3.6000 98.4000 ;
	    RECT 2.8000 83.6000 3.6000 84.4000 ;
	    RECT 12.4000 84.2000 13.2000 97.8000 ;
	    RECT 14.0000 84.2000 14.8000 97.8000 ;
	    RECT 15.6000 84.2000 16.4000 97.8000 ;
	    RECT 17.2000 86.2000 18.0000 97.8000 ;
	    RECT 18.8000 95.6000 19.6000 96.4000 ;
	    RECT 2.9000 68.4000 3.5000 83.6000 ;
	    RECT 2.8000 67.6000 3.6000 68.4000 ;
	    RECT 2.8000 63.6000 3.6000 64.4000 ;
	    RECT 12.4000 64.2000 13.2000 77.8000 ;
	    RECT 14.0000 64.2000 14.8000 77.8000 ;
	    RECT 15.6000 64.2000 16.4000 77.8000 ;
	    RECT 17.2000 64.2000 18.0000 75.8000 ;
	    RECT 18.9000 66.4000 19.5000 95.6000 ;
	    RECT 20.4000 86.2000 21.2000 97.8000 ;
	    RECT 22.1000 94.4000 22.7000 99.7000 ;
	    RECT 22.0000 93.6000 22.8000 94.4000 ;
	    RECT 23.6000 86.2000 24.4000 97.8000 ;
	    RECT 25.2000 84.2000 26.0000 97.8000 ;
	    RECT 26.8000 84.2000 27.6000 97.8000 ;
	    RECT 28.5000 94.4000 29.1000 111.6000 ;
	    RECT 30.0000 109.6000 30.8000 110.4000 ;
	    RECT 30.1000 106.4000 30.7000 109.6000 ;
	    RECT 31.7000 108.4000 32.3000 121.6000 ;
	    RECT 46.1000 110.4000 46.7000 131.6000 ;
	    RECT 58.8000 129.6000 59.6000 130.4000 ;
	    RECT 58.9000 128.4000 59.5000 129.6000 ;
	    RECT 58.8000 127.6000 59.6000 128.4000 ;
	    RECT 54.0000 123.6000 54.8000 124.4000 ;
	    RECT 36.4000 109.6000 37.2000 110.4000 ;
	    RECT 46.0000 109.6000 46.8000 110.4000 ;
	    RECT 31.6000 107.6000 32.4000 108.4000 ;
	    RECT 37.8000 107.6000 38.8000 108.4000 ;
	    RECT 30.0000 105.6000 30.8000 106.4000 ;
	    RECT 34.8000 105.6000 35.6000 106.4000 ;
	    RECT 34.9000 104.4000 35.5000 105.6000 ;
	    RECT 34.8000 103.6000 35.6000 104.4000 ;
	    RECT 38.1000 98.4000 38.7000 107.6000 ;
	    RECT 44.4000 105.6000 45.2000 106.4000 ;
	    RECT 41.2000 103.6000 42.0000 104.4000 ;
	    RECT 41.3000 98.4000 41.9000 103.6000 ;
	    RECT 38.0000 97.6000 38.8000 98.4000 ;
	    RECT 41.2000 97.6000 42.0000 98.4000 ;
	    RECT 39.6000 95.6000 40.4000 96.4000 ;
	    RECT 28.4000 93.6000 29.2000 94.4000 ;
	    RECT 39.7000 92.4000 40.3000 95.6000 ;
	    RECT 41.2000 93.6000 42.0000 94.4000 ;
	    RECT 30.0000 91.6000 30.8000 92.4000 ;
	    RECT 39.6000 91.6000 40.4000 92.4000 ;
	    RECT 18.8000 65.6000 19.6000 66.4000 ;
	    RECT 2.9000 56.3000 3.5000 63.6000 ;
	    RECT 18.9000 58.4000 19.5000 65.6000 ;
	    RECT 20.4000 64.2000 21.2000 75.8000 ;
	    RECT 22.0000 67.6000 22.8000 68.4000 ;
	    RECT 22.1000 62.4000 22.7000 67.6000 ;
	    RECT 23.6000 64.2000 24.4000 75.8000 ;
	    RECT 25.2000 64.2000 26.0000 77.8000 ;
	    RECT 26.8000 64.2000 27.6000 77.8000 ;
	    RECT 30.1000 70.4000 30.7000 91.6000 ;
	    RECT 41.3000 90.4000 41.9000 93.6000 ;
	    RECT 44.5000 92.4000 45.1000 105.6000 ;
	    RECT 47.6000 104.2000 48.4000 117.8000 ;
	    RECT 49.2000 104.2000 50.0000 117.8000 ;
	    RECT 50.8000 104.2000 51.6000 117.8000 ;
	    RECT 52.4000 104.2000 53.2000 115.8000 ;
	    RECT 54.1000 106.4000 54.7000 123.6000 ;
	    RECT 54.0000 105.6000 54.8000 106.4000 ;
	    RECT 55.6000 104.2000 56.4000 115.8000 ;
	    RECT 57.2000 109.6000 58.0000 110.4000 ;
	    RECT 57.3000 108.4000 57.9000 109.6000 ;
	    RECT 57.2000 107.6000 58.0000 108.4000 ;
	    RECT 58.8000 104.2000 59.6000 115.8000 ;
	    RECT 60.4000 104.2000 61.2000 117.8000 ;
	    RECT 62.0000 104.2000 62.8000 117.8000 ;
	    RECT 66.8000 109.6000 67.6000 110.4000 ;
	    RECT 47.6000 97.6000 48.4000 98.4000 ;
	    RECT 70.1000 98.3000 70.7000 131.6000 ;
	    RECT 74.8000 123.6000 75.6000 124.4000 ;
	    RECT 71.6000 105.6000 72.4000 106.4000 ;
	    RECT 68.5000 97.7000 70.7000 98.3000 ;
	    RECT 47.7000 94.4000 48.3000 97.6000 ;
	    RECT 49.2000 95.0000 50.0000 95.8000 ;
	    RECT 50.6000 95.0000 54.8000 95.6000 ;
	    RECT 55.8000 95.0000 56.6000 95.8000 ;
	    RECT 46.0000 93.6000 46.8000 94.4000 ;
	    RECT 47.6000 93.6000 48.4000 94.4000 ;
	    RECT 49.2000 94.2000 49.8000 95.0000 ;
	    RECT 50.6000 94.8000 51.4000 95.0000 ;
	    RECT 54.0000 94.8000 54.8000 95.0000 ;
	    RECT 49.2000 93.6000 54.0000 94.2000 ;
	    RECT 44.4000 91.6000 45.2000 92.4000 ;
	    RECT 46.0000 91.6000 46.8000 92.4000 ;
	    RECT 41.2000 89.6000 42.0000 90.4000 ;
	    RECT 41.3000 74.4000 41.9000 89.6000 ;
	    RECT 41.2000 73.6000 42.0000 74.4000 ;
	    RECT 42.8000 73.6000 43.6000 74.4000 ;
	    RECT 42.9000 72.4000 43.5000 73.6000 ;
	    RECT 42.8000 71.6000 43.6000 72.4000 ;
	    RECT 46.1000 70.4000 46.7000 91.6000 ;
	    RECT 49.2000 90.2000 49.8000 93.6000 ;
	    RECT 53.2000 93.4000 54.0000 93.6000 ;
	    RECT 56.0000 90.2000 56.6000 95.0000 ;
	    RECT 57.2000 93.6000 58.0000 94.4000 ;
	    RECT 58.8000 93.6000 59.6000 94.4000 ;
	    RECT 58.9000 92.4000 59.5000 93.6000 ;
	    RECT 68.5000 92.4000 69.1000 97.7000 ;
	    RECT 70.0000 96.3000 70.8000 96.4000 ;
	    RECT 71.7000 96.3000 72.3000 105.6000 ;
	    RECT 70.0000 95.7000 72.3000 96.3000 ;
	    RECT 70.0000 95.6000 70.8000 95.7000 ;
	    RECT 70.1000 94.4000 70.7000 95.6000 ;
	    RECT 74.9000 94.4000 75.5000 123.6000 ;
	    RECT 76.5000 106.4000 77.1000 141.7000 ;
	    RECT 84.4000 141.6000 85.2000 142.4000 ;
	    RECT 84.5000 138.4000 85.1000 141.6000 ;
	    RECT 84.4000 137.6000 85.2000 138.4000 ;
	    RECT 78.0000 133.6000 78.8000 134.4000 ;
	    RECT 79.6000 133.6000 80.4000 134.4000 ;
	    RECT 81.2000 133.6000 82.0000 134.4000 ;
	    RECT 78.1000 132.4000 78.7000 133.6000 ;
	    RECT 79.7000 132.4000 80.3000 133.6000 ;
	    RECT 81.3000 132.4000 81.9000 133.6000 ;
	    RECT 78.0000 131.6000 78.8000 132.4000 ;
	    RECT 79.6000 131.6000 80.4000 132.4000 ;
	    RECT 81.2000 131.6000 82.0000 132.4000 ;
	    RECT 82.8000 131.6000 83.6000 132.4000 ;
	    RECT 78.1000 118.4000 78.7000 131.6000 ;
	    RECT 78.0000 117.6000 78.8000 118.4000 ;
	    RECT 79.7000 114.4000 80.3000 131.6000 ;
	    RECT 87.7000 128.4000 88.3000 169.6000 ;
	    RECT 87.6000 127.6000 88.4000 128.4000 ;
	    RECT 79.6000 113.6000 80.4000 114.4000 ;
	    RECT 79.6000 107.6000 80.4000 108.4000 ;
	    RECT 79.7000 106.4000 80.3000 107.6000 ;
	    RECT 76.4000 105.6000 77.2000 106.4000 ;
	    RECT 79.6000 105.6000 80.4000 106.4000 ;
	    RECT 90.9000 102.4000 91.5000 173.6000 ;
	    RECT 95.7000 154.4000 96.3000 189.6000 ;
	    RECT 100.5000 186.4000 101.1000 189.6000 ;
	    RECT 105.2000 187.6000 106.0000 188.4000 ;
	    RECT 108.4000 187.6000 109.2000 188.4000 ;
	    RECT 100.4000 185.6000 101.2000 186.4000 ;
	    RECT 105.3000 182.4000 105.9000 187.6000 ;
	    RECT 105.2000 181.6000 106.0000 182.4000 ;
	    RECT 97.2000 179.6000 98.0000 180.4000 ;
	    RECT 105.2000 179.6000 106.0000 180.4000 ;
	    RECT 97.3000 172.4000 97.9000 179.6000 ;
	    RECT 97.2000 171.6000 98.0000 172.4000 ;
	    RECT 95.6000 153.6000 96.4000 154.4000 ;
	    RECT 97.3000 150.4000 97.9000 171.6000 ;
	    RECT 98.8000 164.2000 99.6000 177.8000 ;
	    RECT 100.4000 164.2000 101.2000 177.8000 ;
	    RECT 102.0000 164.2000 102.8000 177.8000 ;
	    RECT 103.6000 166.2000 104.4000 177.8000 ;
	    RECT 105.3000 176.4000 105.9000 179.6000 ;
	    RECT 105.2000 175.6000 106.0000 176.4000 ;
	    RECT 105.3000 162.4000 105.9000 175.6000 ;
	    RECT 106.8000 166.2000 107.6000 177.8000 ;
	    RECT 108.5000 174.4000 109.1000 187.6000 ;
	    RECT 110.1000 182.4000 110.7000 189.6000 ;
	    RECT 113.2000 187.6000 114.0000 188.4000 ;
	    RECT 113.3000 186.4000 113.9000 187.6000 ;
	    RECT 113.2000 185.6000 114.0000 186.4000 ;
	    RECT 110.0000 181.6000 110.8000 182.4000 ;
	    RECT 108.4000 173.6000 109.2000 174.4000 ;
	    RECT 110.0000 166.2000 110.8000 177.8000 ;
	    RECT 111.6000 164.2000 112.4000 177.8000 ;
	    RECT 113.2000 164.2000 114.0000 177.8000 ;
	    RECT 118.1000 172.4000 118.7000 189.6000 ;
	    RECT 122.8000 184.2000 123.6000 197.8000 ;
	    RECT 124.4000 184.2000 125.2000 197.8000 ;
	    RECT 126.0000 184.2000 126.8000 195.8000 ;
	    RECT 127.6000 187.6000 128.4000 188.4000 ;
	    RECT 127.7000 178.4000 128.3000 187.6000 ;
	    RECT 129.2000 184.2000 130.0000 195.8000 ;
	    RECT 130.8000 185.6000 131.6000 186.4000 ;
	    RECT 130.9000 180.4000 131.5000 185.6000 ;
	    RECT 132.4000 184.2000 133.2000 195.8000 ;
	    RECT 134.0000 184.2000 134.8000 197.8000 ;
	    RECT 135.6000 184.2000 136.4000 197.8000 ;
	    RECT 137.2000 184.2000 138.0000 197.8000 ;
	    RECT 153.2000 193.6000 154.0000 194.4000 ;
	    RECT 145.2000 191.6000 146.0000 192.4000 ;
	    RECT 150.0000 191.6000 150.8000 192.4000 ;
	    RECT 134.0000 181.6000 134.8000 182.4000 ;
	    RECT 130.8000 179.6000 131.6000 180.4000 ;
	    RECT 127.6000 177.6000 128.4000 178.4000 ;
	    RECT 130.8000 177.6000 131.6000 178.4000 ;
	    RECT 122.8000 173.6000 123.6000 174.4000 ;
	    RECT 122.9000 172.4000 123.5000 173.6000 ;
	    RECT 134.1000 172.4000 134.7000 181.6000 ;
	    RECT 142.0000 177.6000 142.8000 178.4000 ;
	    RECT 142.1000 176.4000 142.7000 177.6000 ;
	    RECT 142.0000 175.6000 142.8000 176.4000 ;
	    RECT 143.6000 175.6000 144.4000 176.4000 ;
	    RECT 118.0000 171.6000 118.8000 172.4000 ;
	    RECT 122.8000 171.6000 123.6000 172.4000 ;
	    RECT 126.0000 171.6000 126.8000 172.4000 ;
	    RECT 127.6000 171.6000 128.4000 172.4000 ;
	    RECT 129.2000 171.6000 130.0000 172.4000 ;
	    RECT 134.0000 171.6000 134.8000 172.4000 ;
	    RECT 135.6000 171.6000 136.4000 172.4000 ;
	    RECT 138.8000 171.6000 139.6000 172.4000 ;
	    RECT 126.1000 170.4000 126.7000 171.6000 ;
	    RECT 126.0000 169.6000 126.8000 170.4000 ;
	    RECT 129.3000 168.4000 129.9000 171.6000 ;
	    RECT 129.2000 167.6000 130.0000 168.4000 ;
	    RECT 105.2000 161.6000 106.0000 162.4000 ;
	    RECT 113.2000 161.6000 114.0000 162.4000 ;
	    RECT 97.2000 149.6000 98.0000 150.4000 ;
	    RECT 100.4000 149.6000 101.2000 150.4000 ;
	    RECT 95.6000 145.6000 96.4000 146.4000 ;
	    RECT 94.0000 144.3000 94.8000 144.4000 ;
	    RECT 92.5000 143.7000 94.8000 144.3000 ;
	    RECT 92.5000 136.4000 93.1000 143.7000 ;
	    RECT 94.0000 143.6000 94.8000 143.7000 ;
	    RECT 95.7000 138.4000 96.3000 145.6000 ;
	    RECT 95.6000 137.6000 96.4000 138.4000 ;
	    RECT 92.4000 135.6000 93.2000 136.4000 ;
	    RECT 100.5000 132.4000 101.1000 149.6000 ;
	    RECT 105.2000 144.2000 106.0000 157.8000 ;
	    RECT 106.8000 144.2000 107.6000 157.8000 ;
	    RECT 108.4000 144.2000 109.2000 155.8000 ;
	    RECT 110.0000 147.6000 110.8000 148.4000 ;
	    RECT 110.0000 145.6000 110.8000 146.4000 ;
	    RECT 100.4000 131.6000 101.2000 132.4000 ;
	    RECT 100.5000 110.4000 101.1000 131.6000 ;
	    RECT 98.8000 109.6000 99.6000 110.4000 ;
	    RECT 100.4000 109.6000 101.2000 110.4000 ;
	    RECT 78.0000 101.6000 78.8000 102.4000 ;
	    RECT 90.8000 101.6000 91.6000 102.4000 ;
	    RECT 70.0000 93.6000 70.8000 94.4000 ;
	    RECT 74.8000 93.6000 75.6000 94.4000 ;
	    RECT 58.8000 91.6000 59.6000 92.4000 ;
	    RECT 68.4000 91.6000 69.2000 92.4000 ;
	    RECT 49.2000 89.4000 50.0000 90.2000 ;
	    RECT 55.8000 89.4000 56.6000 90.2000 ;
	    RECT 50.8000 83.6000 51.6000 84.4000 ;
	    RECT 68.5000 84.3000 69.1000 91.6000 ;
	    RECT 68.5000 83.7000 70.7000 84.3000 ;
	    RECT 30.0000 69.6000 30.8000 70.4000 ;
	    RECT 31.6000 70.3000 32.4000 70.4000 ;
	    RECT 31.6000 69.7000 33.9000 70.3000 ;
	    RECT 31.6000 69.6000 32.4000 69.7000 ;
	    RECT 22.0000 61.6000 22.8000 62.4000 ;
	    RECT 26.8000 61.6000 27.6000 62.4000 ;
	    RECT 28.4000 61.6000 29.2000 62.4000 ;
	    RECT 22.0000 59.6000 22.8000 60.4000 ;
	    RECT 18.8000 57.6000 19.6000 58.4000 ;
	    RECT 22.1000 56.4000 22.7000 59.6000 ;
	    RECT 26.9000 58.4000 27.5000 61.6000 ;
	    RECT 26.8000 57.6000 27.6000 58.4000 ;
	    RECT 28.5000 56.4000 29.1000 61.6000 ;
	    RECT 4.4000 56.3000 5.2000 56.4000 ;
	    RECT 2.9000 55.7000 5.2000 56.3000 ;
	    RECT 4.4000 55.6000 5.2000 55.7000 ;
	    RECT 22.0000 55.6000 22.8000 56.4000 ;
	    RECT 28.4000 55.6000 29.2000 56.4000 ;
	    RECT 31.6000 55.6000 32.4000 56.4000 ;
	    RECT 4.5000 52.4000 5.1000 55.6000 ;
	    RECT 31.7000 54.4000 32.3000 55.6000 ;
	    RECT 9.2000 53.6000 10.0000 54.4000 ;
	    RECT 31.6000 53.6000 32.4000 54.4000 ;
	    RECT 9.3000 52.4000 9.9000 53.6000 ;
	    RECT 2.8000 51.6000 3.6000 52.4000 ;
	    RECT 4.4000 51.6000 5.2000 52.4000 ;
	    RECT 9.2000 51.6000 10.0000 52.4000 ;
	    RECT 12.4000 51.6000 13.2000 52.4000 ;
	    RECT 17.2000 51.6000 18.0000 52.4000 ;
	    RECT 18.8000 51.6000 19.6000 52.4000 ;
	    RECT 23.6000 51.6000 24.4000 52.4000 ;
	    RECT 30.0000 51.6000 30.8000 52.4000 ;
	    RECT 2.9000 38.4000 3.5000 51.6000 ;
	    RECT 9.3000 38.4000 9.9000 51.6000 ;
	    RECT 17.3000 50.4000 17.9000 51.6000 ;
	    RECT 17.2000 49.6000 18.0000 50.4000 ;
	    RECT 20.4000 49.6000 21.2000 50.4000 ;
	    RECT 23.7000 48.4000 24.3000 51.6000 ;
	    RECT 30.1000 48.4000 30.7000 51.6000 ;
	    RECT 23.6000 47.6000 24.4000 48.4000 ;
	    RECT 30.0000 47.6000 30.8000 48.4000 ;
	    RECT 14.0000 43.6000 14.8000 44.4000 ;
	    RECT 2.8000 37.6000 3.6000 38.4000 ;
	    RECT 6.0000 37.6000 6.8000 38.4000 ;
	    RECT 9.2000 37.6000 10.0000 38.4000 ;
	    RECT 1.2000 25.6000 2.0000 26.4000 ;
	    RECT 1.3000 18.4000 1.9000 25.6000 ;
	    RECT 1.2000 17.6000 2.0000 18.4000 ;
	    RECT 7.6000 17.6000 8.4000 18.4000 ;
	    RECT 14.1000 14.4000 14.7000 43.6000 ;
	    RECT 25.2000 39.6000 26.0000 40.4000 ;
	    RECT 15.6000 24.2000 16.4000 37.8000 ;
	    RECT 17.2000 24.2000 18.0000 37.8000 ;
	    RECT 18.8000 24.2000 19.6000 37.8000 ;
	    RECT 20.4000 24.2000 21.2000 35.8000 ;
	    RECT 22.0000 31.6000 22.8000 32.4000 ;
	    RECT 22.1000 26.4000 22.7000 31.6000 ;
	    RECT 22.0000 25.6000 22.8000 26.4000 ;
	    RECT 22.1000 20.3000 22.7000 25.6000 ;
	    RECT 23.6000 24.2000 24.4000 35.8000 ;
	    RECT 25.3000 28.4000 25.9000 39.6000 ;
	    RECT 25.2000 27.6000 26.0000 28.4000 ;
	    RECT 26.8000 24.2000 27.6000 35.8000 ;
	    RECT 28.4000 24.2000 29.2000 37.8000 ;
	    RECT 30.0000 24.2000 30.8000 37.8000 ;
	    RECT 33.3000 30.4000 33.9000 69.7000 ;
	    RECT 38.0000 69.6000 38.8000 70.4000 ;
	    RECT 46.0000 69.6000 46.8000 70.4000 ;
	    RECT 49.2000 69.6000 50.0000 70.4000 ;
	    RECT 50.9000 68.4000 51.5000 83.6000 ;
	    RECT 68.4000 78.3000 69.2000 78.4000 ;
	    RECT 70.1000 78.3000 70.7000 83.7000 ;
	    RECT 68.4000 77.7000 70.7000 78.3000 ;
	    RECT 68.4000 77.6000 69.2000 77.7000 ;
	    RECT 74.8000 73.6000 75.6000 74.4000 ;
	    RECT 74.9000 72.4000 75.5000 73.6000 ;
	    RECT 54.0000 71.6000 54.8000 72.4000 ;
	    RECT 66.8000 71.6000 67.6000 72.4000 ;
	    RECT 70.0000 71.6000 70.8000 72.4000 ;
	    RECT 74.8000 72.3000 75.6000 72.4000 ;
	    RECT 74.8000 71.7000 77.1000 72.3000 ;
	    RECT 74.8000 71.6000 75.6000 71.7000 ;
	    RECT 55.6000 69.6000 56.4000 70.4000 ;
	    RECT 57.2000 69.6000 58.0000 70.4000 ;
	    RECT 55.7000 68.4000 56.3000 69.6000 ;
	    RECT 57.3000 68.4000 57.9000 69.6000 ;
	    RECT 36.4000 67.6000 37.2000 68.4000 ;
	    RECT 47.6000 68.3000 48.4000 68.4000 ;
	    RECT 47.6000 67.7000 49.9000 68.3000 ;
	    RECT 47.6000 67.6000 48.4000 67.7000 ;
	    RECT 36.5000 60.4000 37.1000 67.6000 ;
	    RECT 41.2000 63.6000 42.0000 64.4000 ;
	    RECT 42.8000 63.6000 43.6000 64.4000 ;
	    RECT 46.0000 63.6000 46.8000 64.4000 ;
	    RECT 36.4000 59.6000 37.2000 60.4000 ;
	    RECT 41.3000 58.4000 41.9000 63.6000 ;
	    RECT 42.9000 62.4000 43.5000 63.6000 ;
	    RECT 42.8000 61.6000 43.6000 62.4000 ;
	    RECT 46.1000 58.4000 46.7000 63.6000 ;
	    RECT 34.8000 57.6000 35.6000 58.4000 ;
	    RECT 41.2000 57.6000 42.0000 58.4000 ;
	    RECT 46.0000 57.6000 46.8000 58.4000 ;
	    RECT 34.9000 56.4000 35.5000 57.6000 ;
	    RECT 34.8000 55.6000 35.6000 56.4000 ;
	    RECT 36.4000 55.6000 37.2000 56.4000 ;
	    RECT 41.2000 55.0000 42.0000 55.8000 ;
	    RECT 42.6000 55.0000 46.8000 55.6000 ;
	    RECT 47.8000 55.0000 48.6000 55.8000 ;
	    RECT 38.0000 53.6000 38.8000 54.4000 ;
	    RECT 41.2000 54.2000 41.8000 55.0000 ;
	    RECT 42.6000 54.8000 43.4000 55.0000 ;
	    RECT 46.0000 54.8000 46.8000 55.0000 ;
	    RECT 41.2000 53.6000 46.0000 54.2000 ;
	    RECT 41.2000 50.2000 41.8000 53.6000 ;
	    RECT 45.2000 53.4000 46.0000 53.6000 ;
	    RECT 48.0000 50.2000 48.6000 55.0000 ;
	    RECT 49.3000 54.4000 49.9000 67.7000 ;
	    RECT 50.8000 67.6000 51.6000 68.4000 ;
	    RECT 55.6000 67.6000 56.4000 68.4000 ;
	    RECT 57.2000 67.6000 58.0000 68.4000 ;
	    RECT 58.8000 67.6000 59.6000 68.4000 ;
	    RECT 54.0000 65.6000 54.8000 66.4000 ;
	    RECT 55.7000 64.4000 56.3000 67.6000 ;
	    RECT 58.9000 66.4000 59.5000 67.6000 ;
	    RECT 66.9000 66.4000 67.5000 71.6000 ;
	    RECT 70.1000 70.4000 70.7000 71.6000 ;
	    RECT 70.0000 69.6000 70.8000 70.4000 ;
	    RECT 73.2000 67.6000 74.0000 68.4000 ;
	    RECT 58.8000 65.6000 59.6000 66.4000 ;
	    RECT 66.8000 65.6000 67.6000 66.4000 ;
	    RECT 55.6000 63.6000 56.4000 64.4000 ;
	    RECT 68.4000 63.6000 69.2000 64.4000 ;
	    RECT 74.8000 63.6000 75.6000 64.4000 ;
	    RECT 52.4000 55.6000 53.2000 56.4000 ;
	    RECT 49.2000 53.6000 50.0000 54.4000 ;
	    RECT 52.5000 52.4000 53.1000 55.6000 ;
	    RECT 68.5000 52.4000 69.1000 63.6000 ;
	    RECT 74.9000 58.4000 75.5000 63.6000 ;
	    RECT 74.8000 57.6000 75.6000 58.4000 ;
	    RECT 71.6000 55.6000 72.4000 56.4000 ;
	    RECT 50.8000 51.6000 51.6000 52.4000 ;
	    RECT 52.4000 51.6000 53.2000 52.4000 ;
	    RECT 57.2000 51.6000 58.0000 52.4000 ;
	    RECT 68.4000 51.6000 69.2000 52.4000 ;
	    RECT 70.0000 51.6000 70.8000 52.4000 ;
	    RECT 41.2000 49.4000 42.0000 50.2000 ;
	    RECT 47.8000 49.4000 48.6000 50.2000 ;
	    RECT 60.4000 47.6000 61.2000 48.4000 ;
	    RECT 34.8000 43.6000 35.6000 44.4000 ;
	    RECT 55.6000 43.6000 56.4000 44.4000 ;
	    RECT 34.9000 40.4000 35.5000 43.6000 ;
	    RECT 34.8000 39.6000 35.6000 40.4000 ;
	    RECT 33.2000 29.6000 34.0000 30.4000 ;
	    RECT 34.8000 29.6000 35.6000 30.4000 ;
	    RECT 44.4000 29.6000 45.2000 30.4000 ;
	    RECT 22.1000 19.7000 24.3000 20.3000 ;
	    RECT 14.0000 13.6000 14.8000 14.4000 ;
	    RECT 17.2000 4.2000 18.0000 17.8000 ;
	    RECT 18.8000 4.2000 19.6000 17.8000 ;
	    RECT 20.4000 4.2000 21.2000 17.8000 ;
	    RECT 22.0000 6.2000 22.8000 17.8000 ;
	    RECT 23.7000 16.4000 24.3000 19.7000 ;
	    RECT 23.6000 15.6000 24.4000 16.4000 ;
	    RECT 25.2000 6.2000 26.0000 17.8000 ;
	    RECT 26.8000 13.6000 27.6000 14.4000 ;
	    RECT 28.4000 6.2000 29.2000 17.8000 ;
	    RECT 30.0000 4.2000 30.8000 17.8000 ;
	    RECT 31.6000 4.2000 32.4000 17.8000 ;
	    RECT 34.9000 12.4000 35.5000 29.6000 ;
	    RECT 44.5000 12.4000 45.1000 29.6000 ;
	    RECT 47.6000 24.2000 48.4000 37.8000 ;
	    RECT 49.2000 24.2000 50.0000 37.8000 ;
	    RECT 50.8000 24.2000 51.6000 35.8000 ;
	    RECT 52.4000 27.6000 53.2000 28.4000 ;
	    RECT 54.0000 24.2000 54.8000 35.8000 ;
	    RECT 55.7000 34.4000 56.3000 43.6000 ;
	    RECT 55.6000 33.6000 56.4000 34.4000 ;
	    RECT 55.6000 31.6000 56.4000 32.4000 ;
	    RECT 55.7000 26.4000 56.3000 31.6000 ;
	    RECT 55.6000 25.6000 56.4000 26.4000 ;
	    RECT 55.7000 20.3000 56.3000 25.6000 ;
	    RECT 57.2000 24.2000 58.0000 35.8000 ;
	    RECT 58.8000 24.2000 59.6000 37.8000 ;
	    RECT 60.4000 24.2000 61.2000 37.8000 ;
	    RECT 62.0000 24.2000 62.8000 37.8000 ;
	    RECT 71.7000 36.3000 72.3000 55.6000 ;
	    RECT 74.8000 43.6000 75.6000 44.4000 ;
	    RECT 71.7000 35.7000 73.9000 36.3000 ;
	    RECT 71.6000 33.6000 72.4000 34.4000 ;
	    RECT 63.6000 29.6000 64.4000 30.4000 ;
	    RECT 55.7000 19.7000 57.9000 20.3000 ;
	    RECT 34.8000 11.6000 35.6000 12.4000 ;
	    RECT 36.4000 11.6000 37.2000 12.4000 ;
	    RECT 44.4000 11.6000 45.2000 12.4000 ;
	    RECT 49.2000 4.2000 50.0000 17.8000 ;
	    RECT 50.8000 4.2000 51.6000 17.8000 ;
	    RECT 52.4000 6.2000 53.2000 17.8000 ;
	    RECT 54.0000 13.6000 54.8000 14.4000 ;
	    RECT 55.6000 6.2000 56.4000 17.8000 ;
	    RECT 57.3000 16.4000 57.9000 19.7000 ;
	    RECT 73.3000 18.4000 73.9000 35.7000 ;
	    RECT 74.9000 32.4000 75.5000 43.6000 ;
	    RECT 76.5000 32.4000 77.1000 71.7000 ;
	    RECT 78.1000 70.4000 78.7000 101.6000 ;
	    RECT 98.9000 98.4000 99.5000 109.6000 ;
	    RECT 102.0000 104.2000 102.8000 117.8000 ;
	    RECT 103.6000 104.2000 104.4000 117.8000 ;
	    RECT 105.2000 104.2000 106.0000 115.8000 ;
	    RECT 106.8000 107.6000 107.6000 108.4000 ;
	    RECT 79.6000 84.2000 80.4000 97.8000 ;
	    RECT 81.2000 84.2000 82.0000 97.8000 ;
	    RECT 82.8000 84.2000 83.6000 97.8000 ;
	    RECT 84.4000 86.2000 85.2000 97.8000 ;
	    RECT 86.0000 95.6000 86.8000 96.4000 ;
	    RECT 87.6000 86.2000 88.4000 97.8000 ;
	    RECT 89.2000 93.6000 90.0000 94.4000 ;
	    RECT 90.8000 86.2000 91.6000 97.8000 ;
	    RECT 92.4000 84.2000 93.2000 97.8000 ;
	    RECT 94.0000 84.2000 94.8000 97.8000 ;
	    RECT 98.8000 97.6000 99.6000 98.4000 ;
	    RECT 98.9000 92.4000 99.5000 97.6000 ;
	    RECT 106.9000 96.3000 107.5000 107.6000 ;
	    RECT 108.4000 104.2000 109.2000 115.8000 ;
	    RECT 110.1000 106.4000 110.7000 145.6000 ;
	    RECT 111.6000 144.2000 112.4000 155.8000 ;
	    RECT 113.3000 146.4000 113.9000 161.6000 ;
	    RECT 113.2000 145.6000 114.0000 146.4000 ;
	    RECT 114.8000 144.2000 115.6000 155.8000 ;
	    RECT 116.4000 144.2000 117.2000 157.8000 ;
	    RECT 118.0000 144.2000 118.8000 157.8000 ;
	    RECT 119.6000 144.2000 120.4000 157.8000 ;
	    RECT 132.4000 151.6000 133.2000 152.4000 ;
	    RECT 129.2000 149.6000 130.2000 150.4000 ;
	    RECT 130.8000 147.6000 131.6000 148.4000 ;
	    RECT 124.4000 145.6000 125.2000 146.4000 ;
	    RECT 111.6000 131.6000 112.4000 132.4000 ;
	    RECT 116.4000 124.2000 117.2000 137.8000 ;
	    RECT 118.0000 124.2000 118.8000 137.8000 ;
	    RECT 119.6000 126.2000 120.4000 137.8000 ;
	    RECT 121.2000 133.6000 122.0000 134.4000 ;
	    RECT 121.3000 124.4000 121.9000 133.6000 ;
	    RECT 122.8000 126.2000 123.6000 137.8000 ;
	    RECT 124.5000 136.4000 125.1000 145.6000 ;
	    RECT 124.4000 135.6000 125.2000 136.4000 ;
	    RECT 126.0000 126.2000 126.8000 137.8000 ;
	    RECT 121.2000 123.6000 122.0000 124.4000 ;
	    RECT 126.0000 123.6000 126.8000 124.4000 ;
	    RECT 127.6000 124.2000 128.4000 137.8000 ;
	    RECT 129.2000 124.2000 130.0000 137.8000 ;
	    RECT 130.8000 124.2000 131.6000 137.8000 ;
	    RECT 126.1000 118.4000 126.7000 123.6000 ;
	    RECT 134.1000 118.4000 134.7000 171.6000 ;
	    RECT 137.2000 169.6000 138.0000 170.4000 ;
	    RECT 145.3000 170.3000 145.9000 191.6000 ;
	    RECT 148.4000 189.6000 149.2000 190.4000 ;
	    RECT 151.6000 189.6000 152.4000 190.4000 ;
	    RECT 146.8000 183.6000 147.6000 184.4000 ;
	    RECT 146.9000 178.4000 147.5000 183.6000 ;
	    RECT 146.8000 177.6000 147.6000 178.4000 ;
	    RECT 143.7000 169.7000 145.9000 170.3000 ;
	    RECT 140.4000 151.6000 141.2000 152.4000 ;
	    RECT 135.6000 149.6000 136.4000 150.4000 ;
	    RECT 140.4000 149.6000 141.2000 150.4000 ;
	    RECT 135.7000 148.4000 136.3000 149.6000 ;
	    RECT 135.6000 147.6000 136.4000 148.4000 ;
	    RECT 140.5000 146.4000 141.1000 149.6000 ;
	    RECT 143.7000 146.4000 144.3000 169.7000 ;
	    RECT 145.2000 163.6000 146.0000 164.4000 ;
	    RECT 145.3000 148.4000 145.9000 163.6000 ;
	    RECT 146.8000 149.6000 147.6000 150.4000 ;
	    RECT 145.2000 147.6000 146.0000 148.4000 ;
	    RECT 146.8000 147.6000 147.6000 148.4000 ;
	    RECT 140.4000 145.6000 141.2000 146.4000 ;
	    RECT 143.6000 145.6000 144.4000 146.4000 ;
	    RECT 143.7000 138.3000 144.3000 145.6000 ;
	    RECT 146.9000 138.4000 147.5000 147.6000 ;
	    RECT 142.1000 137.7000 144.3000 138.3000 ;
	    RECT 142.1000 136.4000 142.7000 137.7000 ;
	    RECT 146.8000 137.6000 147.6000 138.4000 ;
	    RECT 142.0000 135.6000 142.8000 136.4000 ;
	    RECT 143.6000 135.6000 144.4000 136.4000 ;
	    RECT 143.7000 124.4000 144.3000 135.6000 ;
	    RECT 143.6000 123.6000 144.4000 124.4000 ;
	    RECT 110.0000 105.6000 110.8000 106.4000 ;
	    RECT 108.4000 97.6000 109.2000 98.4000 ;
	    RECT 110.1000 96.4000 110.7000 105.6000 ;
	    RECT 111.6000 104.2000 112.4000 115.8000 ;
	    RECT 113.2000 104.2000 114.0000 117.8000 ;
	    RECT 114.8000 104.2000 115.6000 117.8000 ;
	    RECT 116.4000 104.2000 117.2000 117.8000 ;
	    RECT 124.4000 117.6000 125.2000 118.4000 ;
	    RECT 126.0000 117.6000 126.8000 118.4000 ;
	    RECT 134.0000 117.6000 134.8000 118.4000 ;
	    RECT 143.6000 117.6000 144.4000 118.4000 ;
	    RECT 106.9000 95.7000 109.1000 96.3000 ;
	    RECT 106.8000 93.6000 107.6000 94.4000 ;
	    RECT 106.9000 92.4000 107.5000 93.6000 ;
	    RECT 98.8000 91.6000 99.6000 92.4000 ;
	    RECT 106.8000 91.6000 107.6000 92.4000 ;
	    RECT 103.6000 83.6000 104.4000 84.4000 ;
	    RECT 103.7000 80.3000 104.3000 83.6000 ;
	    RECT 108.5000 80.4000 109.1000 95.7000 ;
	    RECT 110.0000 95.6000 110.8000 96.4000 ;
	    RECT 113.2000 93.6000 114.0000 94.4000 ;
	    RECT 113.3000 92.4000 113.9000 93.6000 ;
	    RECT 113.2000 91.6000 114.0000 92.4000 ;
	    RECT 121.2000 91.6000 122.0000 92.4000 ;
	    RECT 124.5000 90.4000 125.1000 117.6000 ;
	    RECT 130.8000 115.6000 131.6000 116.4000 ;
	    RECT 146.8000 115.6000 147.6000 116.4000 ;
	    RECT 130.9000 110.4000 131.5000 115.6000 ;
	    RECT 132.4000 113.6000 133.2000 114.4000 ;
	    RECT 146.9000 112.4000 147.5000 115.6000 ;
	    RECT 148.5000 114.4000 149.1000 189.6000 ;
	    RECT 153.3000 186.4000 153.9000 193.6000 ;
	    RECT 164.4000 189.6000 165.2000 190.4000 ;
	    RECT 150.0000 185.6000 150.8000 186.4000 ;
	    RECT 153.2000 185.6000 154.0000 186.4000 ;
	    RECT 150.1000 148.4000 150.7000 185.6000 ;
	    RECT 151.6000 183.6000 152.4000 184.4000 ;
	    RECT 159.6000 184.3000 160.4000 184.4000 ;
	    RECT 159.6000 183.7000 161.9000 184.3000 ;
	    RECT 159.6000 183.6000 160.4000 183.7000 ;
	    RECT 151.7000 176.4000 152.3000 183.6000 ;
	    RECT 151.6000 175.6000 152.4000 176.4000 ;
	    RECT 158.0000 175.6000 158.8000 176.4000 ;
	    RECT 159.6000 171.6000 160.4000 172.4000 ;
	    RECT 151.6000 169.6000 152.4000 170.4000 ;
	    RECT 151.7000 150.4000 152.3000 169.6000 ;
	    RECT 159.7000 158.4000 160.3000 171.6000 ;
	    RECT 159.6000 157.6000 160.4000 158.4000 ;
	    RECT 161.3000 150.4000 161.9000 183.7000 ;
	    RECT 164.5000 178.4000 165.1000 189.6000 ;
	    RECT 167.6000 183.6000 168.4000 184.4000 ;
	    RECT 177.2000 184.2000 178.0000 197.8000 ;
	    RECT 178.8000 184.2000 179.6000 197.8000 ;
	    RECT 180.4000 184.2000 181.2000 197.8000 ;
	    RECT 182.0000 184.2000 182.8000 195.8000 ;
	    RECT 183.6000 185.6000 184.4000 186.4000 ;
	    RECT 167.7000 180.4000 168.3000 183.6000 ;
	    RECT 167.6000 179.6000 168.4000 180.4000 ;
	    RECT 177.2000 179.6000 178.0000 180.4000 ;
	    RECT 164.4000 177.6000 165.2000 178.4000 ;
	    RECT 166.0000 171.6000 166.8000 172.4000 ;
	    RECT 167.6000 164.2000 168.4000 177.8000 ;
	    RECT 169.2000 164.2000 170.0000 177.8000 ;
	    RECT 170.8000 164.2000 171.6000 177.8000 ;
	    RECT 172.4000 166.2000 173.2000 177.8000 ;
	    RECT 174.0000 175.6000 174.8000 176.4000 ;
	    RECT 174.1000 150.4000 174.7000 175.6000 ;
	    RECT 175.6000 166.2000 176.4000 177.8000 ;
	    RECT 177.3000 174.4000 177.9000 179.6000 ;
	    RECT 177.2000 173.6000 178.0000 174.4000 ;
	    RECT 178.8000 166.2000 179.6000 177.8000 ;
	    RECT 180.4000 164.2000 181.2000 177.8000 ;
	    RECT 182.0000 164.2000 182.8000 177.8000 ;
	    RECT 183.7000 176.4000 184.3000 185.6000 ;
	    RECT 185.2000 184.2000 186.0000 195.8000 ;
	    RECT 188.4000 184.2000 189.2000 195.8000 ;
	    RECT 190.0000 184.2000 190.8000 197.8000 ;
	    RECT 191.6000 184.2000 192.4000 197.8000 ;
	    RECT 194.8000 189.6000 195.6000 190.4000 ;
	    RECT 204.4000 189.6000 205.2000 190.4000 ;
	    RECT 214.0000 189.6000 214.8000 190.4000 ;
	    RECT 218.8000 189.6000 219.6000 190.4000 ;
	    RECT 223.6000 189.6000 224.4000 190.4000 ;
	    RECT 183.6000 175.6000 184.4000 176.4000 ;
	    RECT 194.9000 172.4000 195.5000 189.6000 ;
	    RECT 204.4000 187.6000 205.2000 188.4000 ;
	    RECT 209.2000 187.6000 210.0000 188.4000 ;
	    RECT 188.4000 171.6000 189.2000 172.4000 ;
	    RECT 194.8000 171.6000 195.6000 172.4000 ;
	    RECT 188.5000 150.4000 189.1000 171.6000 ;
	    RECT 199.6000 164.2000 200.4000 177.8000 ;
	    RECT 201.2000 164.2000 202.0000 177.8000 ;
	    RECT 202.8000 166.2000 203.6000 177.8000 ;
	    RECT 204.5000 174.4000 205.1000 187.6000 ;
	    RECT 214.1000 186.4000 214.7000 189.6000 ;
	    RECT 214.0000 185.6000 214.8000 186.4000 ;
	    RECT 220.4000 183.6000 221.2000 184.4000 ;
	    RECT 204.4000 173.6000 205.2000 174.4000 ;
	    RECT 206.0000 166.2000 206.8000 177.8000 ;
	    RECT 207.6000 175.6000 208.4000 176.4000 ;
	    RECT 209.2000 166.2000 210.0000 177.8000 ;
	    RECT 210.8000 164.2000 211.6000 177.8000 ;
	    RECT 212.4000 164.2000 213.2000 177.8000 ;
	    RECT 214.0000 164.2000 214.8000 177.8000 ;
	    RECT 151.6000 149.6000 152.4000 150.4000 ;
	    RECT 161.2000 149.6000 162.0000 150.4000 ;
	    RECT 174.0000 149.6000 174.8000 150.4000 ;
	    RECT 175.6000 149.6000 176.4000 150.4000 ;
	    RECT 180.4000 149.6000 181.2000 150.4000 ;
	    RECT 188.4000 149.6000 189.2000 150.4000 ;
	    RECT 190.0000 149.6000 190.8000 150.4000 ;
	    RECT 150.0000 147.6000 150.8000 148.4000 ;
	    RECT 150.0000 143.6000 150.8000 144.4000 ;
	    RECT 150.1000 134.4000 150.7000 143.6000 ;
	    RECT 174.1000 140.4000 174.7000 149.6000 ;
	    RECT 177.2000 147.6000 178.0000 148.4000 ;
	    RECT 180.4000 147.6000 181.2000 148.4000 ;
	    RECT 180.4000 145.6000 181.2000 146.4000 ;
	    RECT 183.6000 145.6000 184.4000 146.4000 ;
	    RECT 180.5000 144.4000 181.1000 145.6000 ;
	    RECT 180.4000 143.6000 181.2000 144.4000 ;
	    RECT 183.6000 143.6000 184.4000 144.4000 ;
	    RECT 167.6000 139.6000 168.4000 140.4000 ;
	    RECT 174.0000 139.6000 174.8000 140.4000 ;
	    RECT 150.0000 133.6000 150.8000 134.4000 ;
	    RECT 158.0000 131.6000 158.8000 132.4000 ;
	    RECT 158.1000 130.8000 158.7000 131.6000 ;
	    RECT 158.0000 130.0000 158.8000 130.8000 ;
	    RECT 159.6000 124.2000 160.4000 137.8000 ;
	    RECT 161.2000 124.2000 162.0000 137.8000 ;
	    RECT 162.8000 126.2000 163.6000 137.8000 ;
	    RECT 164.4000 133.6000 165.2000 134.4000 ;
	    RECT 166.0000 126.2000 166.8000 137.8000 ;
	    RECT 167.7000 136.4000 168.3000 139.6000 ;
	    RECT 183.7000 138.4000 184.3000 143.6000 ;
	    RECT 167.6000 135.6000 168.4000 136.4000 ;
	    RECT 169.2000 126.2000 170.0000 137.8000 ;
	    RECT 170.8000 124.2000 171.6000 137.8000 ;
	    RECT 172.4000 124.2000 173.2000 137.8000 ;
	    RECT 174.0000 124.2000 174.8000 137.8000 ;
	    RECT 183.6000 137.6000 184.4000 138.4000 ;
	    RECT 190.1000 132.4000 190.7000 149.6000 ;
	    RECT 193.2000 144.2000 194.0000 157.8000 ;
	    RECT 194.8000 144.2000 195.6000 157.8000 ;
	    RECT 196.4000 144.2000 197.2000 155.8000 ;
	    RECT 198.0000 149.6000 198.8000 150.4000 ;
	    RECT 198.1000 148.4000 198.7000 149.6000 ;
	    RECT 198.0000 147.6000 198.8000 148.4000 ;
	    RECT 199.6000 144.2000 200.4000 155.8000 ;
	    RECT 201.2000 145.6000 202.0000 146.4000 ;
	    RECT 201.3000 140.4000 201.9000 145.6000 ;
	    RECT 202.8000 144.2000 203.6000 155.8000 ;
	    RECT 204.4000 144.2000 205.2000 157.8000 ;
	    RECT 206.0000 144.2000 206.8000 157.8000 ;
	    RECT 207.6000 144.2000 208.4000 157.8000 ;
	    RECT 217.2000 145.6000 218.0000 146.4000 ;
	    RECT 201.2000 140.3000 202.0000 140.4000 ;
	    RECT 201.2000 139.7000 203.5000 140.3000 ;
	    RECT 201.2000 139.6000 202.0000 139.7000 ;
	    RECT 190.0000 131.6000 190.8000 132.4000 ;
	    RECT 185.2000 127.6000 186.0000 128.4000 ;
	    RECT 164.4000 117.6000 165.2000 118.4000 ;
	    RECT 148.4000 113.6000 149.2000 114.4000 ;
	    RECT 150.0000 113.6000 150.8000 114.4000 ;
	    RECT 140.4000 111.6000 141.2000 112.4000 ;
	    RECT 145.2000 111.6000 146.0000 112.4000 ;
	    RECT 146.8000 111.6000 147.6000 112.4000 ;
	    RECT 127.6000 109.6000 128.4000 110.4000 ;
	    RECT 130.8000 109.6000 131.6000 110.4000 ;
	    RECT 138.8000 109.6000 139.6000 110.4000 ;
	    RECT 142.0000 109.6000 142.8000 110.4000 ;
	    RECT 126.0000 91.6000 126.8000 92.4000 ;
	    RECT 116.4000 89.6000 117.2000 90.4000 ;
	    RECT 124.4000 89.6000 125.2000 90.4000 ;
	    RECT 116.5000 88.4000 117.1000 89.6000 ;
	    RECT 127.7000 88.4000 128.3000 109.6000 ;
	    RECT 145.3000 106.4000 145.9000 111.6000 ;
	    RECT 150.0000 109.6000 150.8000 110.4000 ;
	    RECT 156.4000 109.6000 157.2000 110.4000 ;
	    RECT 132.4000 105.6000 133.2000 106.4000 ;
	    RECT 135.6000 105.6000 136.4000 106.4000 ;
	    RECT 138.8000 105.6000 139.6000 106.4000 ;
	    RECT 145.2000 105.6000 146.0000 106.4000 ;
	    RECT 153.2000 105.6000 154.0000 106.4000 ;
	    RECT 132.5000 96.4000 133.1000 105.6000 ;
	    RECT 135.7000 104.4000 136.3000 105.6000 ;
	    RECT 135.6000 103.6000 136.4000 104.4000 ;
	    RECT 135.6000 99.6000 136.4000 100.4000 ;
	    RECT 135.7000 98.4000 136.3000 99.6000 ;
	    RECT 135.6000 97.6000 136.4000 98.4000 ;
	    RECT 132.4000 95.6000 133.2000 96.4000 ;
	    RECT 130.8000 91.6000 131.6000 92.4000 ;
	    RECT 116.4000 87.6000 117.2000 88.4000 ;
	    RECT 119.6000 87.6000 120.4000 88.4000 ;
	    RECT 127.6000 87.6000 128.4000 88.4000 ;
	    RECT 118.0000 83.6000 118.8000 84.4000 ;
	    RECT 118.1000 82.4000 118.7000 83.6000 ;
	    RECT 118.0000 81.6000 118.8000 82.4000 ;
	    RECT 103.7000 79.7000 105.9000 80.3000 ;
	    RECT 78.0000 69.6000 78.8000 70.4000 ;
	    RECT 82.8000 69.6000 83.6000 70.4000 ;
	    RECT 79.6000 67.6000 80.4000 68.4000 ;
	    RECT 79.7000 66.4000 80.3000 67.6000 ;
	    RECT 79.6000 65.6000 80.4000 66.4000 ;
	    RECT 79.7000 34.4000 80.3000 65.6000 ;
	    RECT 79.6000 33.6000 80.4000 34.4000 ;
	    RECT 74.8000 31.6000 75.6000 32.4000 ;
	    RECT 76.4000 31.6000 77.2000 32.4000 ;
	    RECT 79.6000 31.6000 80.4000 32.4000 ;
	    RECT 79.7000 28.4000 80.3000 31.6000 ;
	    RECT 82.9000 30.4000 83.5000 69.6000 ;
	    RECT 89.2000 64.2000 90.0000 77.8000 ;
	    RECT 90.8000 64.2000 91.6000 77.8000 ;
	    RECT 92.4000 64.2000 93.2000 75.8000 ;
	    RECT 94.0000 67.6000 94.8000 68.4000 ;
	    RECT 95.6000 64.2000 96.4000 75.8000 ;
	    RECT 97.2000 65.6000 98.0000 66.4000 ;
	    RECT 97.3000 64.4000 97.9000 65.6000 ;
	    RECT 97.2000 63.6000 98.0000 64.4000 ;
	    RECT 98.8000 64.2000 99.6000 75.8000 ;
	    RECT 100.4000 64.2000 101.2000 77.8000 ;
	    RECT 102.0000 64.2000 102.8000 77.8000 ;
	    RECT 103.6000 64.2000 104.4000 77.8000 ;
	    RECT 105.3000 70.4000 105.9000 79.7000 ;
	    RECT 108.4000 79.6000 109.2000 80.4000 ;
	    RECT 118.0000 79.6000 118.8000 80.4000 ;
	    RECT 118.1000 78.4000 118.7000 79.6000 ;
	    RECT 119.7000 78.4000 120.3000 87.6000 ;
	    RECT 126.0000 83.6000 126.8000 84.4000 ;
	    RECT 118.0000 77.6000 118.8000 78.4000 ;
	    RECT 119.6000 77.6000 120.4000 78.4000 ;
	    RECT 105.2000 69.6000 106.0000 70.4000 ;
	    RECT 113.2000 69.6000 114.2000 70.4000 ;
	    RECT 122.8000 69.6000 123.6000 70.4000 ;
	    RECT 126.1000 70.3000 126.7000 83.6000 ;
	    RECT 126.1000 69.7000 128.3000 70.3000 ;
	    RECT 121.2000 67.6000 122.0000 68.4000 ;
	    RECT 121.3000 66.4000 121.9000 67.6000 ;
	    RECT 116.4000 65.6000 117.2000 66.4000 ;
	    RECT 121.2000 65.6000 122.0000 66.4000 ;
	    RECT 103.6000 61.6000 104.4000 62.4000 ;
	    RECT 103.7000 58.4000 104.3000 61.6000 ;
	    RECT 103.6000 57.6000 104.4000 58.4000 ;
	    RECT 102.0000 55.6000 102.8000 56.4000 ;
	    RECT 100.4000 53.6000 101.2000 54.4000 ;
	    RECT 110.0000 53.6000 110.8000 54.4000 ;
	    RECT 106.8000 49.6000 107.6000 50.4000 ;
	    RECT 90.8000 47.6000 91.6000 48.4000 ;
	    RECT 84.4000 33.6000 85.2000 34.4000 ;
	    RECT 82.8000 29.6000 83.6000 30.4000 ;
	    RECT 90.9000 28.4000 91.5000 47.6000 ;
	    RECT 103.6000 43.6000 104.4000 44.4000 ;
	    RECT 100.4000 41.6000 101.2000 42.4000 ;
	    RECT 100.5000 36.4000 101.1000 41.6000 ;
	    RECT 100.4000 35.6000 101.2000 36.4000 ;
	    RECT 92.4000 33.6000 93.2000 34.4000 ;
	    RECT 92.5000 30.4000 93.1000 33.6000 ;
	    RECT 100.5000 32.4000 101.1000 35.6000 ;
	    RECT 103.7000 34.4000 104.3000 43.6000 ;
	    RECT 105.2000 35.6000 106.0000 36.4000 ;
	    RECT 108.4000 35.6000 109.2000 36.4000 ;
	    RECT 108.5000 34.4000 109.1000 35.6000 ;
	    RECT 103.6000 33.6000 104.4000 34.4000 ;
	    RECT 108.4000 33.6000 109.2000 34.4000 ;
	    RECT 97.2000 31.6000 98.0000 32.4000 ;
	    RECT 100.4000 31.6000 101.2000 32.4000 ;
	    RECT 110.1000 32.3000 110.7000 53.6000 ;
	    RECT 111.6000 51.6000 112.4000 52.4000 ;
	    RECT 113.2000 51.6000 114.0000 52.4000 ;
	    RECT 111.7000 50.4000 112.3000 51.6000 ;
	    RECT 113.3000 50.4000 113.9000 51.6000 ;
	    RECT 111.6000 49.6000 112.4000 50.4000 ;
	    RECT 113.2000 49.6000 114.0000 50.4000 ;
	    RECT 114.8000 47.6000 115.6000 48.4000 ;
	    RECT 113.2000 43.6000 114.0000 44.4000 ;
	    RECT 113.3000 34.4000 113.9000 43.6000 ;
	    RECT 116.5000 36.4000 117.1000 65.6000 ;
	    RECT 121.2000 51.6000 122.0000 52.4000 ;
	    RECT 121.3000 50.4000 121.9000 51.6000 ;
	    RECT 122.9000 50.4000 123.5000 69.6000 ;
	    RECT 127.7000 68.4000 128.3000 69.7000 ;
	    RECT 129.2000 69.6000 130.0000 70.4000 ;
	    RECT 129.3000 68.4000 129.9000 69.6000 ;
	    RECT 132.5000 68.4000 133.1000 95.6000 ;
	    RECT 138.9000 92.4000 139.5000 105.6000 ;
	    RECT 145.3000 100.4000 145.9000 105.6000 ;
	    RECT 156.5000 104.4000 157.1000 109.6000 ;
	    RECT 164.5000 108.4000 165.1000 117.6000 ;
	    RECT 183.6000 115.6000 184.4000 116.4000 ;
	    RECT 174.0000 111.6000 174.8000 112.4000 ;
	    RECT 185.3000 110.4000 185.9000 127.6000 ;
	    RECT 194.8000 124.2000 195.6000 137.8000 ;
	    RECT 196.4000 124.2000 197.2000 137.8000 ;
	    RECT 198.0000 126.2000 198.8000 137.8000 ;
	    RECT 199.6000 133.6000 200.4000 134.4000 ;
	    RECT 199.7000 122.4000 200.3000 133.6000 ;
	    RECT 201.2000 126.2000 202.0000 137.8000 ;
	    RECT 202.9000 136.4000 203.5000 139.7000 ;
	    RECT 202.8000 135.6000 203.6000 136.4000 ;
	    RECT 204.4000 126.2000 205.2000 137.8000 ;
	    RECT 206.0000 124.2000 206.8000 137.8000 ;
	    RECT 207.6000 124.2000 208.4000 137.8000 ;
	    RECT 209.2000 124.2000 210.0000 137.8000 ;
	    RECT 218.8000 123.6000 219.6000 124.4000 ;
	    RECT 194.8000 121.6000 195.6000 122.4000 ;
	    RECT 199.6000 121.6000 200.4000 122.4000 ;
	    RECT 194.9000 118.4000 195.5000 121.6000 ;
	    RECT 194.8000 117.6000 195.6000 118.4000 ;
	    RECT 191.6000 113.6000 192.4000 114.4000 ;
	    RECT 191.7000 112.4000 192.3000 113.6000 ;
	    RECT 186.8000 111.6000 187.6000 112.4000 ;
	    RECT 191.6000 111.6000 192.4000 112.4000 ;
	    RECT 198.0000 111.6000 198.8000 112.4000 ;
	    RECT 186.9000 110.4000 187.5000 111.6000 ;
	    RECT 198.1000 110.4000 198.7000 111.6000 ;
	    RECT 218.9000 110.4000 219.5000 123.6000 ;
	    RECT 170.8000 109.6000 171.6000 110.4000 ;
	    RECT 182.0000 109.6000 182.8000 110.4000 ;
	    RECT 185.2000 109.6000 186.0000 110.4000 ;
	    RECT 186.8000 109.6000 187.6000 110.4000 ;
	    RECT 198.0000 109.6000 198.8000 110.4000 ;
	    RECT 209.2000 109.6000 210.0000 110.4000 ;
	    RECT 218.8000 109.6000 219.6000 110.4000 ;
	    RECT 164.4000 107.6000 165.2000 108.4000 ;
	    RECT 169.2000 107.6000 170.0000 108.4000 ;
	    RECT 167.6000 105.6000 168.4000 106.4000 ;
	    RECT 170.9000 106.3000 171.5000 109.6000 ;
	    RECT 175.6000 107.6000 176.4000 108.4000 ;
	    RECT 180.4000 107.6000 181.2000 108.4000 ;
	    RECT 170.9000 105.7000 173.1000 106.3000 ;
	    RECT 156.4000 103.6000 157.2000 104.4000 ;
	    RECT 166.0000 103.6000 166.8000 104.4000 ;
	    RECT 145.2000 99.6000 146.0000 100.4000 ;
	    RECT 138.8000 91.6000 139.6000 92.4000 ;
	    RECT 143.6000 91.6000 144.4000 92.4000 ;
	    RECT 143.7000 90.4000 144.3000 91.6000 ;
	    RECT 143.6000 89.6000 144.4000 90.4000 ;
	    RECT 135.6000 83.6000 136.4000 84.4000 ;
	    RECT 145.2000 84.2000 146.0000 97.8000 ;
	    RECT 146.8000 84.2000 147.6000 97.8000 ;
	    RECT 148.4000 84.2000 149.2000 97.8000 ;
	    RECT 150.0000 86.2000 150.8000 97.8000 ;
	    RECT 151.6000 95.6000 152.4000 96.4000 ;
	    RECT 151.7000 84.3000 152.3000 95.6000 ;
	    RECT 153.2000 86.2000 154.0000 97.8000 ;
	    RECT 154.8000 93.6000 155.6000 94.4000 ;
	    RECT 156.4000 86.2000 157.2000 97.8000 ;
	    RECT 151.7000 83.7000 153.9000 84.3000 ;
	    RECT 158.0000 84.2000 158.8000 97.8000 ;
	    RECT 159.6000 84.2000 160.4000 97.8000 ;
	    RECT 161.2000 91.6000 162.0000 92.4000 ;
	    RECT 124.4000 67.6000 125.2000 68.4000 ;
	    RECT 126.0000 67.6000 126.8000 68.4000 ;
	    RECT 127.6000 67.6000 128.4000 68.4000 ;
	    RECT 129.2000 67.6000 130.0000 68.4000 ;
	    RECT 132.4000 67.6000 133.2000 68.4000 ;
	    RECT 124.5000 62.4000 125.1000 67.6000 ;
	    RECT 124.4000 61.6000 125.2000 62.4000 ;
	    RECT 126.1000 58.4000 126.7000 67.6000 ;
	    RECT 127.6000 63.6000 128.4000 64.4000 ;
	    RECT 126.0000 57.6000 126.8000 58.4000 ;
	    RECT 127.7000 52.4000 128.3000 63.6000 ;
	    RECT 127.6000 51.6000 128.4000 52.4000 ;
	    RECT 119.6000 49.6000 120.4000 50.4000 ;
	    RECT 121.2000 49.6000 122.0000 50.4000 ;
	    RECT 122.8000 49.6000 123.6000 50.4000 ;
	    RECT 119.7000 48.4000 120.3000 49.6000 ;
	    RECT 119.6000 47.6000 120.4000 48.4000 ;
	    RECT 116.4000 35.6000 117.2000 36.4000 ;
	    RECT 113.2000 33.6000 114.0000 34.4000 ;
	    RECT 116.4000 33.6000 117.2000 34.4000 ;
	    RECT 108.5000 31.7000 110.7000 32.3000 ;
	    RECT 92.4000 29.6000 93.2000 30.4000 ;
	    RECT 79.6000 27.6000 80.4000 28.4000 ;
	    RECT 81.2000 27.6000 82.0000 28.4000 ;
	    RECT 89.2000 27.6000 90.0000 28.4000 ;
	    RECT 90.8000 27.6000 91.6000 28.4000 ;
	    RECT 95.6000 27.6000 96.4000 28.4000 ;
	    RECT 89.3000 26.4000 89.9000 27.6000 ;
	    RECT 89.2000 25.6000 90.0000 26.4000 ;
	    RECT 57.2000 15.6000 58.0000 16.4000 ;
	    RECT 58.8000 6.2000 59.6000 17.8000 ;
	    RECT 60.4000 4.2000 61.2000 17.8000 ;
	    RECT 62.0000 4.2000 62.8000 17.8000 ;
	    RECT 63.6000 4.2000 64.4000 17.8000 ;
	    RECT 73.2000 17.6000 74.0000 18.4000 ;
	    RECT 89.3000 12.4000 89.9000 25.6000 ;
	    RECT 90.9000 14.4000 91.5000 27.6000 ;
	    RECT 97.3000 26.4000 97.9000 31.6000 ;
	    RECT 98.8000 29.6000 99.6000 30.4000 ;
	    RECT 102.0000 29.6000 102.8000 30.4000 ;
	    RECT 97.2000 25.6000 98.0000 26.4000 ;
	    RECT 90.8000 13.6000 91.6000 14.4000 ;
	    RECT 89.2000 11.6000 90.0000 12.4000 ;
	    RECT 102.0000 4.2000 102.8000 17.8000 ;
	    RECT 103.6000 4.2000 104.4000 17.8000 ;
	    RECT 105.2000 4.2000 106.0000 17.8000 ;
	    RECT 106.8000 6.2000 107.6000 17.8000 ;
	    RECT 108.5000 16.4000 109.1000 31.7000 ;
	    RECT 111.6000 31.6000 112.4000 32.4000 ;
	    RECT 110.0000 29.6000 110.8000 30.4000 ;
	    RECT 110.1000 28.4000 110.7000 29.6000 ;
	    RECT 111.7000 28.4000 112.3000 31.6000 ;
	    RECT 116.5000 30.4000 117.1000 33.6000 ;
	    RECT 119.7000 30.4000 120.3000 47.6000 ;
	    RECT 121.2000 45.6000 122.0000 46.4000 ;
	    RECT 122.9000 42.4000 123.5000 49.6000 ;
	    RECT 122.8000 41.6000 123.6000 42.4000 ;
	    RECT 116.4000 29.6000 117.2000 30.4000 ;
	    RECT 119.6000 29.6000 120.4000 30.4000 ;
	    RECT 110.0000 27.6000 110.8000 28.4000 ;
	    RECT 111.6000 27.6000 112.4000 28.4000 ;
	    RECT 118.0000 27.6000 118.8000 28.4000 ;
	    RECT 118.1000 26.4000 118.7000 27.6000 ;
	    RECT 110.0000 25.6000 110.8000 26.4000 ;
	    RECT 118.0000 25.6000 118.8000 26.4000 ;
	    RECT 119.6000 25.6000 120.4000 26.4000 ;
	    RECT 113.2000 23.6000 114.0000 24.4000 ;
	    RECT 126.0000 23.6000 126.8000 24.4000 ;
	    RECT 113.3000 20.3000 113.9000 23.6000 ;
	    RECT 111.7000 19.7000 113.9000 20.3000 ;
	    RECT 108.4000 15.6000 109.2000 16.4000 ;
	    RECT 110.0000 6.2000 110.8000 17.8000 ;
	    RECT 111.7000 14.4000 112.3000 19.7000 ;
	    RECT 126.1000 18.4000 126.7000 23.6000 ;
	    RECT 111.6000 13.6000 112.4000 14.4000 ;
	    RECT 113.2000 6.2000 114.0000 17.8000 ;
	    RECT 114.8000 4.2000 115.6000 17.8000 ;
	    RECT 116.4000 4.2000 117.2000 17.8000 ;
	    RECT 126.0000 17.6000 126.8000 18.4000 ;
	    RECT 129.3000 16.4000 129.9000 67.6000 ;
	    RECT 135.7000 66.4000 136.3000 83.6000 ;
	    RECT 151.6000 69.6000 152.4000 70.4000 ;
	    RECT 135.6000 65.6000 136.4000 66.4000 ;
	    RECT 134.0000 63.6000 134.8000 64.4000 ;
	    RECT 142.0000 63.6000 142.8000 64.4000 ;
	    RECT 134.1000 48.4000 134.7000 63.6000 ;
	    RECT 134.0000 47.6000 134.8000 48.4000 ;
	    RECT 135.6000 44.2000 136.4000 57.8000 ;
	    RECT 137.2000 44.2000 138.0000 57.8000 ;
	    RECT 138.8000 44.2000 139.6000 57.8000 ;
	    RECT 140.4000 46.2000 141.2000 57.8000 ;
	    RECT 142.1000 56.4000 142.7000 63.6000 ;
	    RECT 142.0000 55.6000 142.8000 56.4000 ;
	    RECT 142.1000 54.4000 142.7000 55.6000 ;
	    RECT 142.0000 53.6000 142.8000 54.4000 ;
	    RECT 134.0000 29.6000 134.8000 30.4000 ;
	    RECT 130.8000 17.6000 131.6000 18.4000 ;
	    RECT 126.0000 15.6000 126.8000 16.4000 ;
	    RECT 129.2000 15.6000 130.0000 16.4000 ;
	    RECT 126.1000 12.4000 126.7000 15.6000 ;
	    RECT 130.9000 12.4000 131.5000 17.6000 ;
	    RECT 134.1000 12.4000 134.7000 29.6000 ;
	    RECT 135.6000 24.2000 136.4000 37.8000 ;
	    RECT 137.2000 24.2000 138.0000 37.8000 ;
	    RECT 138.8000 24.2000 139.6000 37.8000 ;
	    RECT 140.4000 24.2000 141.2000 35.8000 ;
	    RECT 142.1000 26.4000 142.7000 53.6000 ;
	    RECT 143.6000 46.2000 144.4000 57.8000 ;
	    RECT 145.2000 53.6000 146.0000 54.4000 ;
	    RECT 146.8000 46.2000 147.6000 57.8000 ;
	    RECT 148.4000 44.2000 149.2000 57.8000 ;
	    RECT 150.0000 44.2000 150.8000 57.8000 ;
	    RECT 151.7000 52.4000 152.3000 69.6000 ;
	    RECT 153.3000 64.4000 153.9000 83.7000 ;
	    RECT 153.2000 63.6000 154.0000 64.4000 ;
	    RECT 156.4000 64.2000 157.2000 77.8000 ;
	    RECT 158.0000 64.2000 158.8000 77.8000 ;
	    RECT 159.6000 64.2000 160.4000 75.8000 ;
	    RECT 161.3000 70.4000 161.9000 91.6000 ;
	    RECT 161.2000 69.6000 162.0000 70.4000 ;
	    RECT 161.2000 67.6000 162.0000 68.4000 ;
	    RECT 162.8000 64.2000 163.6000 75.8000 ;
	    RECT 164.4000 65.6000 165.2000 66.4000 ;
	    RECT 164.5000 64.4000 165.1000 65.6000 ;
	    RECT 164.4000 63.6000 165.2000 64.4000 ;
	    RECT 166.0000 64.2000 166.8000 75.8000 ;
	    RECT 167.6000 64.2000 168.4000 77.8000 ;
	    RECT 169.2000 64.2000 170.0000 77.8000 ;
	    RECT 170.8000 64.2000 171.6000 77.8000 ;
	    RECT 164.4000 57.6000 165.2000 58.4000 ;
	    RECT 164.5000 54.4000 165.1000 57.6000 ;
	    RECT 164.4000 53.6000 165.2000 54.4000 ;
	    RECT 167.6000 53.6000 168.4000 54.4000 ;
	    RECT 170.8000 53.6000 171.6000 54.4000 ;
	    RECT 172.5000 52.4000 173.1000 105.7000 ;
	    RECT 175.7000 104.4000 176.3000 107.6000 ;
	    RECT 175.6000 103.6000 176.4000 104.4000 ;
	    RECT 177.2000 103.6000 178.0000 104.4000 ;
	    RECT 177.3000 94.4000 177.9000 103.6000 ;
	    RECT 180.5000 102.4000 181.1000 107.6000 ;
	    RECT 185.3000 106.4000 185.9000 109.6000 ;
	    RECT 196.4000 107.6000 197.2000 108.4000 ;
	    RECT 185.2000 105.6000 186.0000 106.4000 ;
	    RECT 196.5000 104.4000 197.1000 107.6000 ;
	    RECT 196.4000 103.6000 197.2000 104.4000 ;
	    RECT 180.4000 101.6000 181.2000 102.4000 ;
	    RECT 177.2000 93.6000 178.0000 94.4000 ;
	    RECT 177.2000 91.6000 178.0000 92.4000 ;
	    RECT 182.0000 84.2000 182.8000 97.8000 ;
	    RECT 183.6000 84.2000 184.4000 97.8000 ;
	    RECT 185.2000 86.2000 186.0000 97.8000 ;
	    RECT 186.8000 93.6000 187.6000 94.4000 ;
	    RECT 186.9000 84.4000 187.5000 93.6000 ;
	    RECT 188.4000 86.2000 189.2000 97.8000 ;
	    RECT 190.0000 95.6000 190.8000 96.4000 ;
	    RECT 191.6000 86.2000 192.4000 97.8000 ;
	    RECT 186.8000 83.6000 187.6000 84.4000 ;
	    RECT 191.6000 83.6000 192.4000 84.4000 ;
	    RECT 193.2000 84.2000 194.0000 97.8000 ;
	    RECT 194.8000 84.2000 195.6000 97.8000 ;
	    RECT 196.4000 84.2000 197.2000 97.8000 ;
	    RECT 191.7000 78.4000 192.3000 83.6000 ;
	    RECT 191.6000 77.6000 192.4000 78.4000 ;
	    RECT 188.4000 75.6000 189.2000 76.4000 ;
	    RECT 188.5000 72.4000 189.1000 75.6000 ;
	    RECT 194.8000 73.6000 195.6000 74.4000 ;
	    RECT 194.9000 72.4000 195.5000 73.6000 ;
	    RECT 198.1000 72.4000 198.7000 109.6000 ;
	    RECT 218.9000 108.4000 219.5000 109.6000 ;
	    RECT 204.4000 107.6000 205.2000 108.4000 ;
	    RECT 210.8000 107.6000 211.6000 108.4000 ;
	    RECT 218.8000 107.6000 219.6000 108.4000 ;
	    RECT 204.5000 106.4000 205.1000 107.6000 ;
	    RECT 210.9000 106.4000 211.5000 107.6000 ;
	    RECT 204.4000 105.6000 205.2000 106.4000 ;
	    RECT 210.8000 105.6000 211.6000 106.4000 ;
	    RECT 218.8000 105.6000 219.6000 106.4000 ;
	    RECT 207.6000 103.6000 208.4000 104.4000 ;
	    RECT 212.4000 103.6000 213.2000 104.4000 ;
	    RECT 207.7000 92.4000 208.3000 103.6000 ;
	    RECT 209.2000 101.6000 210.0000 102.4000 ;
	    RECT 209.3000 98.4000 209.9000 101.6000 ;
	    RECT 209.2000 97.6000 210.0000 98.4000 ;
	    RECT 212.4000 93.6000 213.2000 94.4000 ;
	    RECT 207.6000 91.6000 208.4000 92.4000 ;
	    RECT 206.0000 83.6000 206.8000 84.4000 ;
	    RECT 206.1000 80.4000 206.7000 83.6000 ;
	    RECT 206.0000 79.6000 206.8000 80.4000 ;
	    RECT 206.0000 73.6000 206.8000 74.4000 ;
	    RECT 185.2000 71.6000 186.0000 72.4000 ;
	    RECT 188.4000 71.6000 189.2000 72.4000 ;
	    RECT 190.0000 71.6000 190.8000 72.4000 ;
	    RECT 194.8000 71.6000 195.6000 72.4000 ;
	    RECT 198.0000 71.6000 198.8000 72.4000 ;
	    RECT 202.8000 71.6000 203.6000 72.4000 ;
	    RECT 175.6000 69.6000 176.4000 70.4000 ;
	    RECT 185.2000 69.6000 186.0000 70.4000 ;
	    RECT 175.7000 58.4000 176.3000 69.6000 ;
	    RECT 190.1000 68.4000 190.7000 71.6000 ;
	    RECT 202.9000 70.4000 203.5000 71.6000 ;
	    RECT 207.7000 70.4000 208.3000 91.6000 ;
	    RECT 209.2000 89.6000 210.0000 90.4000 ;
	    RECT 212.5000 88.4000 213.1000 93.6000 ;
	    RECT 215.6000 91.6000 216.4000 92.4000 ;
	    RECT 217.2000 91.6000 218.0000 92.4000 ;
	    RECT 215.6000 89.6000 216.4000 90.4000 ;
	    RECT 212.4000 87.6000 213.2000 88.4000 ;
	    RECT 217.3000 82.4000 217.9000 91.6000 ;
	    RECT 218.9000 90.3000 219.5000 105.6000 ;
	    RECT 220.5000 94.4000 221.1000 183.6000 ;
	    RECT 223.7000 178.4000 224.3000 189.6000 ;
	    RECT 223.6000 177.6000 224.4000 178.4000 ;
	    RECT 222.0000 109.6000 222.8000 110.4000 ;
	    RECT 220.4000 93.6000 221.2000 94.4000 ;
	    RECT 222.1000 92.4000 222.7000 109.6000 ;
	    RECT 222.0000 91.6000 222.8000 92.4000 ;
	    RECT 220.4000 90.3000 221.2000 90.4000 ;
	    RECT 218.9000 89.7000 221.2000 90.3000 ;
	    RECT 217.2000 81.6000 218.0000 82.4000 ;
	    RECT 210.8000 75.6000 211.6000 76.4000 ;
	    RECT 212.4000 73.6000 213.2000 74.4000 ;
	    RECT 217.2000 73.6000 218.0000 74.4000 ;
	    RECT 209.2000 71.6000 210.0000 72.4000 ;
	    RECT 191.6000 69.6000 192.4000 70.4000 ;
	    RECT 198.0000 69.6000 198.8000 70.4000 ;
	    RECT 201.2000 69.6000 202.0000 70.4000 ;
	    RECT 202.8000 69.6000 203.6000 70.4000 ;
	    RECT 206.0000 69.6000 206.8000 70.4000 ;
	    RECT 207.6000 69.6000 208.4000 70.4000 ;
	    RECT 210.8000 69.6000 211.6000 70.4000 ;
	    RECT 212.4000 69.6000 213.2000 70.4000 ;
	    RECT 217.2000 69.6000 218.0000 70.4000 ;
	    RECT 183.6000 67.6000 184.4000 68.4000 ;
	    RECT 190.0000 67.6000 190.8000 68.4000 ;
	    RECT 185.2000 65.6000 186.0000 66.4000 ;
	    RECT 180.4000 63.6000 181.2000 64.4000 ;
	    RECT 175.6000 57.6000 176.4000 58.4000 ;
	    RECT 177.2000 53.6000 178.0000 54.4000 ;
	    RECT 183.6000 53.6000 184.4000 54.4000 ;
	    RECT 183.7000 52.4000 184.3000 53.6000 ;
	    RECT 151.6000 51.6000 152.4000 52.4000 ;
	    RECT 166.0000 51.6000 166.8000 52.4000 ;
	    RECT 172.4000 51.6000 173.2000 52.4000 ;
	    RECT 177.2000 51.6000 178.0000 52.4000 ;
	    RECT 180.4000 51.6000 181.2000 52.4000 ;
	    RECT 182.0000 51.6000 182.8000 52.4000 ;
	    RECT 183.6000 51.6000 184.4000 52.4000 ;
	    RECT 142.0000 25.6000 142.8000 26.4000 ;
	    RECT 142.1000 24.4000 142.7000 25.6000 ;
	    RECT 142.0000 23.6000 142.8000 24.4000 ;
	    RECT 143.6000 24.2000 144.4000 35.8000 ;
	    RECT 145.2000 27.6000 146.0000 28.4000 ;
	    RECT 135.6000 17.6000 136.4000 18.4000 ;
	    RECT 137.2000 17.6000 138.0000 18.4000 ;
	    RECT 135.7000 16.4000 136.3000 17.6000 ;
	    RECT 145.3000 16.4000 145.9000 27.6000 ;
	    RECT 146.8000 24.2000 147.6000 35.8000 ;
	    RECT 148.4000 24.2000 149.2000 37.8000 ;
	    RECT 150.0000 24.2000 150.8000 37.8000 ;
	    RECT 151.7000 30.4000 152.3000 51.6000 ;
	    RECT 169.2000 49.6000 170.0000 50.4000 ;
	    RECT 169.3000 44.4000 169.9000 49.6000 ;
	    RECT 172.5000 46.4000 173.1000 51.6000 ;
	    RECT 177.3000 50.4000 177.9000 51.6000 ;
	    RECT 177.2000 49.6000 178.0000 50.4000 ;
	    RECT 180.5000 48.4000 181.1000 51.6000 ;
	    RECT 180.4000 47.6000 181.2000 48.4000 ;
	    RECT 172.4000 45.6000 173.2000 46.4000 ;
	    RECT 169.2000 43.6000 170.0000 44.4000 ;
	    RECT 151.6000 29.6000 152.4000 30.4000 ;
	    RECT 172.4000 29.6000 173.2000 30.4000 ;
	    RECT 146.8000 17.6000 147.6000 18.4000 ;
	    RECT 135.6000 15.6000 136.4000 16.4000 ;
	    RECT 145.2000 15.6000 146.0000 16.4000 ;
	    RECT 135.7000 12.4000 136.3000 15.6000 ;
	    RECT 146.9000 14.4000 147.5000 17.6000 ;
	    RECT 140.4000 13.6000 141.2000 14.4000 ;
	    RECT 146.8000 13.6000 147.6000 14.4000 ;
	    RECT 151.7000 12.4000 152.3000 29.6000 ;
	    RECT 161.2000 27.6000 162.0000 28.4000 ;
	    RECT 167.6000 27.6000 168.4000 28.4000 ;
	    RECT 161.3000 20.4000 161.9000 27.6000 ;
	    RECT 162.8000 25.6000 163.6000 26.4000 ;
	    RECT 169.2000 25.6000 170.0000 26.4000 ;
	    RECT 170.8000 25.6000 171.6000 26.4000 ;
	    RECT 161.2000 19.6000 162.0000 20.4000 ;
	    RECT 156.4000 17.6000 157.2000 18.4000 ;
	    RECT 153.2000 15.6000 154.0000 16.4000 ;
	    RECT 156.5000 12.4000 157.1000 17.6000 ;
	    RECT 161.3000 14.4000 161.9000 19.6000 ;
	    RECT 169.3000 16.4000 169.9000 25.6000 ;
	    RECT 169.2000 15.6000 170.0000 16.4000 ;
	    RECT 172.5000 14.4000 173.1000 29.6000 ;
	    RECT 175.6000 27.6000 176.4000 28.4000 ;
	    RECT 177.2000 27.6000 178.0000 28.4000 ;
	    RECT 180.4000 27.6000 181.2000 28.4000 ;
	    RECT 175.7000 26.4000 176.3000 27.6000 ;
	    RECT 175.6000 25.6000 176.4000 26.4000 ;
	    RECT 177.2000 25.6000 178.0000 26.4000 ;
	    RECT 182.1000 22.4000 182.7000 51.6000 ;
	    RECT 183.6000 49.6000 184.4000 50.4000 ;
	    RECT 183.7000 48.4000 184.3000 49.6000 ;
	    RECT 183.6000 47.6000 184.4000 48.4000 ;
	    RECT 185.3000 32.4000 185.9000 65.6000 ;
	    RECT 186.8000 63.6000 187.6000 64.4000 ;
	    RECT 186.9000 56.4000 187.5000 63.6000 ;
	    RECT 190.1000 58.4000 190.7000 67.6000 ;
	    RECT 191.7000 58.4000 192.3000 69.6000 ;
	    RECT 201.3000 66.4000 201.9000 69.6000 ;
	    RECT 206.1000 66.4000 206.7000 69.6000 ;
	    RECT 212.5000 66.4000 213.1000 69.6000 ;
	    RECT 196.4000 65.6000 197.2000 66.4000 ;
	    RECT 201.2000 65.6000 202.0000 66.4000 ;
	    RECT 202.8000 65.6000 203.6000 66.4000 ;
	    RECT 206.0000 65.6000 206.8000 66.4000 ;
	    RECT 212.4000 65.6000 213.2000 66.4000 ;
	    RECT 190.0000 57.6000 190.8000 58.4000 ;
	    RECT 191.6000 57.6000 192.4000 58.4000 ;
	    RECT 199.6000 57.6000 200.4000 58.4000 ;
	    RECT 186.8000 55.6000 187.6000 56.4000 ;
	    RECT 190.2000 55.6000 191.0000 55.8000 ;
	    RECT 186.9000 52.4000 187.5000 55.6000 ;
	    RECT 190.2000 55.0000 195.8000 55.6000 ;
	    RECT 196.4000 55.0000 197.2000 55.8000 ;
	    RECT 188.4000 53.6000 189.2000 54.4000 ;
	    RECT 186.8000 51.6000 187.6000 52.4000 ;
	    RECT 188.5000 48.4000 189.1000 53.6000 ;
	    RECT 190.2000 50.2000 190.8000 55.0000 ;
	    RECT 191.6000 54.8000 192.4000 55.0000 ;
	    RECT 195.0000 54.8000 195.8000 55.0000 ;
	    RECT 196.6000 54.2000 197.2000 55.0000 ;
	    RECT 191.6000 53.6000 197.2000 54.2000 ;
	    RECT 198.0000 53.6000 198.8000 54.4000 ;
	    RECT 191.6000 52.2000 192.2000 53.6000 ;
	    RECT 191.4000 51.4000 192.2000 52.2000 ;
	    RECT 194.8000 51.6000 195.6000 52.4000 ;
	    RECT 190.2000 49.4000 191.0000 50.2000 ;
	    RECT 188.4000 47.6000 189.2000 48.4000 ;
	    RECT 185.2000 31.6000 186.0000 32.4000 ;
	    RECT 182.0000 21.6000 182.8000 22.4000 ;
	    RECT 185.3000 20.4000 185.9000 31.6000 ;
	    RECT 188.5000 26.4000 189.1000 47.6000 ;
	    RECT 194.9000 36.4000 195.5000 51.6000 ;
	    RECT 196.6000 50.2000 197.2000 53.6000 ;
	    RECT 199.7000 50.4000 200.3000 57.6000 ;
	    RECT 202.9000 52.4000 203.5000 65.6000 ;
	    RECT 212.5000 58.4000 213.1000 65.6000 ;
	    RECT 215.6000 63.6000 216.4000 64.4000 ;
	    RECT 212.4000 57.6000 213.2000 58.4000 ;
	    RECT 210.8000 55.6000 211.6000 56.4000 ;
	    RECT 204.4000 53.6000 205.2000 54.4000 ;
	    RECT 214.0000 53.6000 214.8000 54.4000 ;
	    RECT 202.8000 51.6000 203.6000 52.4000 ;
	    RECT 204.4000 51.6000 205.2000 52.4000 ;
	    RECT 196.4000 49.4000 197.2000 50.2000 ;
	    RECT 199.6000 49.6000 200.4000 50.4000 ;
	    RECT 190.0000 35.6000 190.8000 36.4000 ;
	    RECT 193.2000 35.6000 194.0000 36.4000 ;
	    RECT 194.8000 35.6000 195.6000 36.4000 ;
	    RECT 190.1000 28.4000 190.7000 35.6000 ;
	    RECT 193.3000 34.4000 193.9000 35.6000 ;
	    RECT 193.2000 33.6000 194.0000 34.4000 ;
	    RECT 194.8000 33.6000 195.6000 34.4000 ;
	    RECT 191.6000 31.6000 192.4000 32.4000 ;
	    RECT 198.0000 32.3000 198.8000 32.4000 ;
	    RECT 199.7000 32.3000 200.3000 49.6000 ;
	    RECT 210.8000 43.6000 211.6000 44.4000 ;
	    RECT 210.9000 38.4000 211.5000 43.6000 ;
	    RECT 210.8000 37.6000 211.6000 38.4000 ;
	    RECT 215.7000 38.3000 216.3000 63.6000 ;
	    RECT 218.9000 58.4000 219.5000 89.7000 ;
	    RECT 220.4000 89.6000 221.2000 89.7000 ;
	    RECT 222.0000 87.6000 222.8000 88.4000 ;
	    RECT 223.6000 87.6000 224.4000 88.4000 ;
	    RECT 222.1000 86.4000 222.7000 87.6000 ;
	    RECT 222.0000 85.6000 222.8000 86.4000 ;
	    RECT 223.7000 84.3000 224.3000 87.6000 ;
	    RECT 222.1000 83.7000 224.3000 84.3000 ;
	    RECT 222.1000 76.3000 222.7000 83.7000 ;
	    RECT 223.6000 81.6000 224.4000 82.4000 ;
	    RECT 223.7000 78.4000 224.3000 81.6000 ;
	    RECT 223.6000 77.6000 224.4000 78.4000 ;
	    RECT 222.1000 75.7000 224.3000 76.3000 ;
	    RECT 218.8000 57.6000 219.6000 58.4000 ;
	    RECT 217.2000 55.6000 218.0000 56.4000 ;
	    RECT 223.7000 38.4000 224.3000 75.7000 ;
	    RECT 214.1000 37.7000 216.3000 38.3000 ;
	    RECT 214.1000 32.4000 214.7000 37.7000 ;
	    RECT 223.6000 37.6000 224.4000 38.4000 ;
	    RECT 215.6000 35.6000 216.4000 36.4000 ;
	    RECT 215.7000 34.4000 216.3000 35.6000 ;
	    RECT 215.6000 33.6000 216.4000 34.4000 ;
	    RECT 217.2000 33.6000 218.0000 34.4000 ;
	    RECT 198.0000 31.7000 200.3000 32.3000 ;
	    RECT 198.0000 31.6000 198.8000 31.7000 ;
	    RECT 214.0000 31.6000 214.8000 32.4000 ;
	    RECT 217.3000 30.4000 217.9000 33.6000 ;
	    RECT 193.2000 29.6000 194.0000 30.4000 ;
	    RECT 201.2000 29.6000 202.0000 30.4000 ;
	    RECT 206.0000 29.6000 206.8000 30.4000 ;
	    RECT 210.8000 29.6000 211.6000 30.4000 ;
	    RECT 217.2000 29.6000 218.0000 30.4000 ;
	    RECT 190.0000 27.6000 190.8000 28.4000 ;
	    RECT 188.4000 25.6000 189.2000 26.4000 ;
	    RECT 193.3000 24.4000 193.9000 29.6000 ;
	    RECT 199.6000 27.6000 200.4000 28.4000 ;
	    RECT 199.7000 26.4000 200.3000 27.6000 ;
	    RECT 199.6000 25.6000 200.4000 26.4000 ;
	    RECT 204.4000 25.6000 205.2000 26.4000 ;
	    RECT 186.8000 23.6000 187.6000 24.4000 ;
	    RECT 188.4000 23.6000 189.2000 24.4000 ;
	    RECT 193.2000 23.6000 194.0000 24.4000 ;
	    RECT 185.2000 19.6000 186.0000 20.4000 ;
	    RECT 161.2000 13.6000 162.0000 14.4000 ;
	    RECT 172.4000 13.6000 173.2000 14.4000 ;
	    RECT 121.2000 11.6000 122.0000 12.4000 ;
	    RECT 126.0000 11.6000 126.8000 12.4000 ;
	    RECT 130.8000 11.6000 131.6000 12.4000 ;
	    RECT 134.0000 11.6000 134.8000 12.4000 ;
	    RECT 135.6000 11.6000 136.4000 12.4000 ;
	    RECT 142.0000 11.6000 142.8000 12.4000 ;
	    RECT 151.6000 11.6000 152.4000 12.4000 ;
	    RECT 156.4000 11.6000 157.2000 12.4000 ;
	    RECT 161.3000 10.4000 161.9000 13.6000 ;
	    RECT 178.8000 11.6000 179.6000 12.4000 ;
	    RECT 151.6000 9.6000 152.4000 10.4000 ;
	    RECT 161.2000 9.6000 162.0000 10.4000 ;
	    RECT 180.4000 4.2000 181.2000 17.8000 ;
	    RECT 182.0000 4.2000 182.8000 17.8000 ;
	    RECT 183.6000 4.2000 184.4000 17.8000 ;
	    RECT 185.2000 6.2000 186.0000 17.8000 ;
	    RECT 186.9000 16.4000 187.5000 23.6000 ;
	    RECT 188.5000 20.3000 189.1000 23.6000 ;
	    RECT 188.5000 19.7000 190.7000 20.3000 ;
	    RECT 186.8000 15.6000 187.6000 16.4000 ;
	    RECT 188.4000 6.2000 189.2000 17.8000 ;
	    RECT 190.1000 14.4000 190.7000 19.7000 ;
	    RECT 190.0000 13.6000 190.8000 14.4000 ;
	    RECT 191.6000 6.2000 192.4000 17.8000 ;
	    RECT 193.2000 4.2000 194.0000 17.8000 ;
	    RECT 194.8000 4.2000 195.6000 17.8000 ;
	    RECT 206.1000 16.4000 206.7000 29.6000 ;
	    RECT 209.2000 23.6000 210.0000 24.4000 ;
	    RECT 209.3000 18.4000 209.9000 23.6000 ;
	    RECT 217.3000 18.4000 217.9000 29.6000 ;
	    RECT 220.4000 21.6000 221.2000 22.4000 ;
	    RECT 209.2000 17.6000 210.0000 18.4000 ;
	    RECT 210.8000 17.6000 211.6000 18.4000 ;
	    RECT 217.2000 17.6000 218.0000 18.4000 ;
	    RECT 206.0000 15.6000 206.8000 16.4000 ;
	    RECT 218.8000 15.6000 219.6000 16.4000 ;
	    RECT 206.1000 12.4000 206.7000 15.6000 ;
	    RECT 220.5000 12.4000 221.1000 21.6000 ;
	    RECT 206.0000 11.6000 206.8000 12.4000 ;
	    RECT 220.4000 11.6000 221.2000 12.4000 ;
	    RECT 209.2000 9.6000 210.0000 10.4000 ;
	    RECT 212.4000 9.6000 213.2000 10.4000 ;
         LAYER metal3 ;
	    RECT 145.2000 192.3000 146.0000 192.4000 ;
	    RECT 150.0000 192.3000 150.8000 192.4000 ;
	    RECT 145.2000 191.7000 150.8000 192.3000 ;
	    RECT 145.2000 191.6000 146.0000 191.7000 ;
	    RECT 150.0000 191.6000 150.8000 191.7000 ;
	    RECT 89.2000 190.3000 90.0000 190.4000 ;
	    RECT 100.4000 190.3000 101.2000 190.4000 ;
	    RECT 89.2000 189.7000 101.2000 190.3000 ;
	    RECT 89.2000 189.6000 90.0000 189.7000 ;
	    RECT 100.4000 189.6000 101.2000 189.7000 ;
	    RECT 148.4000 190.3000 149.2000 190.4000 ;
	    RECT 151.6000 190.3000 152.4000 190.4000 ;
	    RECT 148.4000 189.7000 152.4000 190.3000 ;
	    RECT 148.4000 189.6000 149.2000 189.7000 ;
	    RECT 151.6000 189.6000 152.4000 189.7000 ;
	    RECT 204.4000 190.3000 205.2000 190.4000 ;
	    RECT 214.0000 190.3000 214.8000 190.4000 ;
	    RECT 218.8000 190.3000 219.6000 190.4000 ;
	    RECT 223.6000 190.3000 224.4000 190.4000 ;
	    RECT 204.4000 189.7000 209.9000 190.3000 ;
	    RECT 204.4000 189.6000 205.2000 189.7000 ;
	    RECT 209.3000 188.4000 209.9000 189.7000 ;
	    RECT 214.0000 189.7000 224.4000 190.3000 ;
	    RECT 214.0000 189.6000 214.8000 189.7000 ;
	    RECT 218.8000 189.6000 219.6000 189.7000 ;
	    RECT 223.6000 189.6000 224.4000 189.7000 ;
	    RECT 14.0000 188.3000 14.8000 188.4000 ;
	    RECT 26.8000 188.3000 27.6000 188.4000 ;
	    RECT 14.0000 187.7000 27.6000 188.3000 ;
	    RECT 14.0000 187.6000 14.8000 187.7000 ;
	    RECT 26.8000 187.6000 27.6000 187.7000 ;
	    RECT 90.8000 188.3000 91.6000 188.4000 ;
	    RECT 113.2000 188.3000 114.0000 188.4000 ;
	    RECT 90.8000 187.7000 114.0000 188.3000 ;
	    RECT 90.8000 187.6000 91.6000 187.7000 ;
	    RECT 113.2000 187.6000 114.0000 187.7000 ;
	    RECT 151.6000 188.3000 152.4000 188.4000 ;
	    RECT 209.2000 188.3000 210.0000 188.4000 ;
	    RECT 151.6000 187.7000 210.0000 188.3000 ;
	    RECT 151.6000 187.6000 152.4000 187.7000 ;
	    RECT 209.2000 187.6000 210.0000 187.7000 ;
	    RECT 150.0000 186.3000 150.8000 186.4000 ;
	    RECT 153.2000 186.3000 154.0000 186.4000 ;
	    RECT 150.0000 185.7000 154.0000 186.3000 ;
	    RECT 150.0000 185.6000 150.8000 185.7000 ;
	    RECT 153.2000 185.6000 154.0000 185.7000 ;
	    RECT 52.4000 184.3000 53.2000 184.4000 ;
	    RECT 57.2000 184.3000 58.0000 184.4000 ;
	    RECT 52.4000 183.7000 58.0000 184.3000 ;
	    RECT 52.4000 183.6000 53.2000 183.7000 ;
	    RECT 57.2000 183.6000 58.0000 183.7000 ;
	    RECT 151.6000 184.3000 152.4000 184.4000 ;
	    RECT 167.6000 184.3000 168.4000 184.4000 ;
	    RECT 151.6000 183.7000 168.4000 184.3000 ;
	    RECT 151.6000 183.6000 152.4000 183.7000 ;
	    RECT 167.6000 183.6000 168.4000 183.7000 ;
	    RECT 17.2000 182.3000 18.0000 182.4000 ;
	    RECT 73.2000 182.3000 74.0000 182.4000 ;
	    RECT 81.2000 182.3000 82.0000 182.4000 ;
	    RECT 105.2000 182.3000 106.0000 182.4000 ;
	    RECT 110.0000 182.3000 110.8000 182.4000 ;
	    RECT 134.0000 182.3000 134.8000 182.4000 ;
	    RECT 151.6000 182.3000 152.4000 182.4000 ;
	    RECT 17.2000 181.7000 152.4000 182.3000 ;
	    RECT 17.2000 181.6000 18.0000 181.7000 ;
	    RECT 73.2000 181.6000 74.0000 181.7000 ;
	    RECT 81.2000 181.6000 82.0000 181.7000 ;
	    RECT 105.2000 181.6000 106.0000 181.7000 ;
	    RECT 110.0000 181.6000 110.8000 181.7000 ;
	    RECT 134.0000 181.6000 134.8000 181.7000 ;
	    RECT 151.6000 181.6000 152.4000 181.7000 ;
	    RECT 36.4000 180.3000 37.2000 180.4000 ;
	    RECT 49.2000 180.3000 50.0000 180.4000 ;
	    RECT 81.2000 180.3000 82.0000 180.4000 ;
	    RECT 97.2000 180.3000 98.0000 180.4000 ;
	    RECT 36.4000 179.7000 98.0000 180.3000 ;
	    RECT 36.4000 179.6000 37.2000 179.7000 ;
	    RECT 49.2000 179.6000 50.0000 179.7000 ;
	    RECT 81.2000 179.6000 82.0000 179.7000 ;
	    RECT 97.2000 179.6000 98.0000 179.7000 ;
	    RECT 105.2000 180.3000 106.0000 180.4000 ;
	    RECT 130.8000 180.3000 131.6000 180.4000 ;
	    RECT 105.2000 179.7000 131.6000 180.3000 ;
	    RECT 105.2000 179.6000 106.0000 179.7000 ;
	    RECT 130.8000 179.6000 131.6000 179.7000 ;
	    RECT 167.6000 180.3000 168.4000 180.4000 ;
	    RECT 177.2000 180.3000 178.0000 180.4000 ;
	    RECT 167.6000 179.7000 178.0000 180.3000 ;
	    RECT 167.6000 179.6000 168.4000 179.7000 ;
	    RECT 177.2000 179.6000 178.0000 179.7000 ;
	    RECT 39.6000 178.3000 40.4000 178.4000 ;
	    RECT 78.0000 178.3000 78.8000 178.4000 ;
	    RECT 39.6000 177.7000 78.8000 178.3000 ;
	    RECT 39.6000 177.6000 40.4000 177.7000 ;
	    RECT 78.0000 177.6000 78.8000 177.7000 ;
	    RECT 127.6000 178.3000 128.4000 178.4000 ;
	    RECT 130.8000 178.3000 131.6000 178.4000 ;
	    RECT 127.6000 177.7000 131.6000 178.3000 ;
	    RECT 127.6000 177.6000 128.4000 177.7000 ;
	    RECT 130.8000 177.6000 131.6000 177.7000 ;
	    RECT 142.0000 178.3000 142.8000 178.4000 ;
	    RECT 146.8000 178.3000 147.6000 178.4000 ;
	    RECT 164.4000 178.3000 165.2000 178.4000 ;
	    RECT 142.0000 177.7000 165.2000 178.3000 ;
	    RECT 142.0000 177.6000 142.8000 177.7000 ;
	    RECT 146.8000 177.6000 147.6000 177.7000 ;
	    RECT 164.4000 177.6000 165.2000 177.7000 ;
	    RECT 23.6000 176.3000 24.4000 176.4000 ;
	    RECT 36.4000 176.3000 37.2000 176.4000 ;
	    RECT 68.4000 176.3000 69.2000 176.4000 ;
	    RECT 23.6000 175.7000 69.2000 176.3000 ;
	    RECT 23.6000 175.6000 24.4000 175.7000 ;
	    RECT 36.4000 175.6000 37.2000 175.7000 ;
	    RECT 68.4000 175.6000 69.2000 175.7000 ;
	    RECT 79.6000 176.3000 80.4000 176.4000 ;
	    RECT 84.4000 176.3000 85.2000 176.4000 ;
	    RECT 79.6000 175.7000 85.2000 176.3000 ;
	    RECT 79.6000 175.6000 80.4000 175.7000 ;
	    RECT 84.4000 175.6000 85.2000 175.7000 ;
	    RECT 143.6000 176.3000 144.4000 176.4000 ;
	    RECT 158.0000 176.3000 158.8000 176.4000 ;
	    RECT 143.6000 175.7000 158.8000 176.3000 ;
	    RECT 143.6000 175.6000 144.4000 175.7000 ;
	    RECT 158.0000 175.6000 158.8000 175.7000 ;
	    RECT 174.0000 176.3000 174.8000 176.4000 ;
	    RECT 183.6000 176.3000 184.4000 176.4000 ;
	    RECT 207.6000 176.3000 208.4000 176.4000 ;
	    RECT 174.0000 175.7000 208.4000 176.3000 ;
	    RECT 174.0000 175.6000 174.8000 175.7000 ;
	    RECT 183.6000 175.6000 184.4000 175.7000 ;
	    RECT 207.6000 175.6000 208.4000 175.7000 ;
	    RECT 76.4000 174.3000 77.2000 174.4000 ;
	    RECT 71.7000 173.7000 77.2000 174.3000 ;
	    RECT 71.7000 172.4000 72.3000 173.7000 ;
	    RECT 76.4000 173.6000 77.2000 173.7000 ;
	    RECT 81.2000 174.3000 82.0000 174.4000 ;
	    RECT 90.8000 174.3000 91.6000 174.4000 ;
	    RECT 81.2000 173.7000 91.6000 174.3000 ;
	    RECT 81.2000 173.6000 82.0000 173.7000 ;
	    RECT 90.8000 173.6000 91.6000 173.7000 ;
	    RECT 57.2000 172.3000 58.0000 172.4000 ;
	    RECT 71.6000 172.3000 72.4000 172.4000 ;
	    RECT 57.2000 171.7000 72.4000 172.3000 ;
	    RECT 57.2000 171.6000 58.0000 171.7000 ;
	    RECT 71.6000 171.6000 72.4000 171.7000 ;
	    RECT 74.8000 172.3000 75.6000 172.4000 ;
	    RECT 82.8000 172.3000 83.6000 172.4000 ;
	    RECT 74.8000 171.7000 83.6000 172.3000 ;
	    RECT 74.8000 171.6000 75.6000 171.7000 ;
	    RECT 82.8000 171.6000 83.6000 171.7000 ;
	    RECT 118.0000 172.3000 118.8000 172.4000 ;
	    RECT 122.8000 172.3000 123.6000 172.4000 ;
	    RECT 118.0000 171.7000 123.6000 172.3000 ;
	    RECT 118.0000 171.6000 118.8000 171.7000 ;
	    RECT 122.8000 171.6000 123.6000 171.7000 ;
	    RECT 127.6000 172.3000 128.4000 172.4000 ;
	    RECT 134.0000 172.3000 134.8000 172.4000 ;
	    RECT 127.6000 171.7000 134.8000 172.3000 ;
	    RECT 127.6000 171.6000 128.4000 171.7000 ;
	    RECT 134.0000 171.6000 134.8000 171.7000 ;
	    RECT 135.6000 172.3000 136.4000 172.4000 ;
	    RECT 138.8000 172.3000 139.6000 172.4000 ;
	    RECT 135.6000 171.7000 139.6000 172.3000 ;
	    RECT 135.6000 171.6000 136.4000 171.7000 ;
	    RECT 138.8000 171.6000 139.6000 171.7000 ;
	    RECT 159.6000 172.3000 160.4000 172.4000 ;
	    RECT 166.0000 172.3000 166.8000 172.4000 ;
	    RECT 159.6000 171.7000 166.8000 172.3000 ;
	    RECT 159.6000 171.6000 160.4000 171.7000 ;
	    RECT 166.0000 171.6000 166.8000 171.7000 ;
	    RECT 188.4000 172.3000 189.2000 172.4000 ;
	    RECT 194.8000 172.3000 195.6000 172.4000 ;
	    RECT 188.4000 171.7000 195.6000 172.3000 ;
	    RECT 188.4000 171.6000 189.2000 171.7000 ;
	    RECT 194.8000 171.6000 195.6000 171.7000 ;
	    RECT 116.4000 170.3000 117.2000 170.4000 ;
	    RECT 126.0000 170.3000 126.8000 170.4000 ;
	    RECT 137.2000 170.3000 138.0000 170.4000 ;
	    RECT 151.6000 170.3000 152.4000 170.4000 ;
	    RECT 116.4000 169.7000 152.4000 170.3000 ;
	    RECT 116.4000 169.6000 117.2000 169.7000 ;
	    RECT 126.0000 169.6000 126.8000 169.7000 ;
	    RECT 137.2000 169.6000 138.0000 169.7000 ;
	    RECT 151.6000 169.6000 152.4000 169.7000 ;
	    RECT 60.4000 168.3000 61.2000 168.4000 ;
	    RECT 129.2000 168.3000 130.0000 168.4000 ;
	    RECT 60.4000 167.7000 130.0000 168.3000 ;
	    RECT 60.4000 167.6000 61.2000 167.7000 ;
	    RECT 129.2000 167.6000 130.0000 167.7000 ;
	    RECT 4.4000 166.3000 5.2000 166.4000 ;
	    RECT 20.4000 166.3000 21.2000 166.4000 ;
	    RECT 54.0000 166.3000 54.8000 166.4000 ;
	    RECT 4.4000 165.7000 54.8000 166.3000 ;
	    RECT 4.4000 165.6000 5.2000 165.7000 ;
	    RECT 20.4000 165.6000 21.2000 165.7000 ;
	    RECT 54.0000 165.6000 54.8000 165.7000 ;
	    RECT 105.2000 162.3000 106.0000 162.4000 ;
	    RECT 113.2000 162.3000 114.0000 162.4000 ;
	    RECT 105.2000 161.7000 114.0000 162.3000 ;
	    RECT 105.2000 161.6000 106.0000 161.7000 ;
	    RECT 113.2000 161.6000 114.0000 161.7000 ;
	    RECT 17.2000 159.6000 18.0000 160.4000 ;
	    RECT 132.4000 152.3000 133.2000 152.4000 ;
	    RECT 140.4000 152.3000 141.2000 152.4000 ;
	    RECT 132.4000 151.7000 141.2000 152.3000 ;
	    RECT 132.4000 151.6000 133.2000 151.7000 ;
	    RECT 140.4000 151.6000 141.2000 151.7000 ;
	    RECT 36.4000 150.3000 37.2000 150.4000 ;
	    RECT 39.6000 150.3000 40.4000 150.4000 ;
	    RECT 36.4000 149.7000 40.4000 150.3000 ;
	    RECT 36.4000 149.6000 37.2000 149.7000 ;
	    RECT 39.6000 149.6000 40.4000 149.7000 ;
	    RECT 44.4000 150.3000 45.2000 150.4000 ;
	    RECT 52.4000 150.3000 53.2000 150.4000 ;
	    RECT 74.8000 150.3000 75.6000 150.4000 ;
	    RECT 44.4000 149.7000 75.6000 150.3000 ;
	    RECT 44.4000 149.6000 45.2000 149.7000 ;
	    RECT 52.4000 149.6000 53.2000 149.7000 ;
	    RECT 74.8000 149.6000 75.6000 149.7000 ;
	    RECT 86.0000 150.3000 86.8000 150.4000 ;
	    RECT 97.2000 150.3000 98.0000 150.4000 ;
	    RECT 86.0000 149.7000 98.0000 150.3000 ;
	    RECT 86.0000 149.6000 86.8000 149.7000 ;
	    RECT 97.2000 149.6000 98.0000 149.7000 ;
	    RECT 129.2000 150.3000 130.0000 150.4000 ;
	    RECT 140.4000 150.3000 141.2000 150.4000 ;
	    RECT 146.8000 150.3000 147.6000 150.4000 ;
	    RECT 129.2000 149.7000 147.6000 150.3000 ;
	    RECT 129.2000 149.6000 130.0000 149.7000 ;
	    RECT 140.4000 149.6000 141.2000 149.7000 ;
	    RECT 146.8000 149.6000 147.6000 149.7000 ;
	    RECT 161.2000 150.3000 162.0000 150.4000 ;
	    RECT 175.6000 150.3000 176.4000 150.4000 ;
	    RECT 161.2000 149.7000 176.4000 150.3000 ;
	    RECT 161.2000 149.6000 162.0000 149.7000 ;
	    RECT 175.6000 149.6000 176.4000 149.7000 ;
	    RECT 180.4000 150.3000 181.2000 150.4000 ;
	    RECT 198.0000 150.3000 198.8000 150.4000 ;
	    RECT 180.4000 149.7000 198.8000 150.3000 ;
	    RECT 180.4000 149.6000 181.2000 149.7000 ;
	    RECT 198.0000 149.6000 198.8000 149.7000 ;
	    RECT 14.0000 148.3000 14.8000 148.4000 ;
	    RECT 26.8000 148.3000 27.6000 148.4000 ;
	    RECT 14.0000 147.7000 27.6000 148.3000 ;
	    RECT 14.0000 147.6000 14.8000 147.7000 ;
	    RECT 26.8000 147.6000 27.6000 147.7000 ;
	    RECT 39.6000 148.3000 40.4000 148.4000 ;
	    RECT 41.2000 148.3000 42.0000 148.4000 ;
	    RECT 39.6000 147.7000 42.0000 148.3000 ;
	    RECT 39.6000 147.6000 40.4000 147.7000 ;
	    RECT 41.2000 147.6000 42.0000 147.7000 ;
	    RECT 46.0000 148.3000 46.8000 148.4000 ;
	    RECT 54.0000 148.3000 54.8000 148.4000 ;
	    RECT 46.0000 147.7000 54.8000 148.3000 ;
	    RECT 46.0000 147.6000 46.8000 147.7000 ;
	    RECT 54.0000 147.6000 54.8000 147.7000 ;
	    RECT 110.0000 148.3000 110.8000 148.4000 ;
	    RECT 130.8000 148.3000 131.6000 148.4000 ;
	    RECT 110.0000 147.7000 131.6000 148.3000 ;
	    RECT 110.0000 147.6000 110.8000 147.7000 ;
	    RECT 130.8000 147.6000 131.6000 147.7000 ;
	    RECT 135.6000 148.3000 136.4000 148.4000 ;
	    RECT 145.2000 148.3000 146.0000 148.4000 ;
	    RECT 135.6000 147.7000 146.0000 148.3000 ;
	    RECT 135.6000 147.6000 136.4000 147.7000 ;
	    RECT 145.2000 147.6000 146.0000 147.7000 ;
	    RECT 146.8000 148.3000 147.6000 148.4000 ;
	    RECT 150.0000 148.3000 150.8000 148.4000 ;
	    RECT 146.8000 147.7000 150.8000 148.3000 ;
	    RECT 146.8000 147.6000 147.6000 147.7000 ;
	    RECT 150.0000 147.6000 150.8000 147.7000 ;
	    RECT 177.2000 148.3000 178.0000 148.4000 ;
	    RECT 180.4000 148.3000 181.2000 148.4000 ;
	    RECT 177.2000 147.7000 181.2000 148.3000 ;
	    RECT 177.2000 147.6000 178.0000 147.7000 ;
	    RECT 180.4000 147.6000 181.2000 147.7000 ;
	    RECT 23.6000 146.3000 24.4000 146.4000 ;
	    RECT 36.4000 146.3000 37.2000 146.4000 ;
	    RECT 23.6000 145.7000 37.2000 146.3000 ;
	    RECT 23.6000 145.6000 24.4000 145.7000 ;
	    RECT 36.4000 145.6000 37.2000 145.7000 ;
	    RECT 42.8000 146.3000 43.6000 146.4000 ;
	    RECT 47.6000 146.3000 48.4000 146.4000 ;
	    RECT 42.8000 145.7000 48.4000 146.3000 ;
	    RECT 42.8000 145.6000 43.6000 145.7000 ;
	    RECT 47.6000 145.6000 48.4000 145.7000 ;
	    RECT 95.6000 146.3000 96.4000 146.4000 ;
	    RECT 110.0000 146.3000 110.8000 146.4000 ;
	    RECT 113.2000 146.3000 114.0000 146.4000 ;
	    RECT 124.4000 146.3000 125.2000 146.4000 ;
	    RECT 95.6000 145.7000 125.2000 146.3000 ;
	    RECT 95.6000 145.6000 96.4000 145.7000 ;
	    RECT 110.0000 145.6000 110.8000 145.7000 ;
	    RECT 113.2000 145.6000 114.0000 145.7000 ;
	    RECT 124.4000 145.6000 125.2000 145.7000 ;
	    RECT 183.6000 146.3000 184.4000 146.4000 ;
	    RECT 217.2000 146.3000 218.0000 146.4000 ;
	    RECT 183.6000 145.7000 218.0000 146.3000 ;
	    RECT 183.6000 145.6000 184.4000 145.7000 ;
	    RECT 217.2000 145.6000 218.0000 145.7000 ;
	    RECT 180.4000 144.3000 181.2000 144.4000 ;
	    RECT 183.6000 144.3000 184.4000 144.4000 ;
	    RECT 180.4000 143.7000 184.4000 144.3000 ;
	    RECT 180.4000 143.6000 181.2000 143.7000 ;
	    RECT 183.6000 143.6000 184.4000 143.7000 ;
	    RECT 74.8000 142.3000 75.6000 142.4000 ;
	    RECT 84.4000 142.3000 85.2000 142.4000 ;
	    RECT 74.8000 141.7000 85.2000 142.3000 ;
	    RECT 74.8000 141.6000 75.6000 141.7000 ;
	    RECT 84.4000 141.6000 85.2000 141.7000 ;
	    RECT 167.6000 140.3000 168.4000 140.4000 ;
	    RECT 174.0000 140.3000 174.8000 140.4000 ;
	    RECT 201.2000 140.3000 202.0000 140.4000 ;
	    RECT 167.6000 139.7000 202.0000 140.3000 ;
	    RECT 167.6000 139.6000 168.4000 139.7000 ;
	    RECT 174.0000 139.6000 174.8000 139.7000 ;
	    RECT 201.2000 139.6000 202.0000 139.7000 ;
	    RECT 4.4000 138.3000 5.2000 138.4000 ;
	    RECT 20.4000 138.3000 21.2000 138.4000 ;
	    RECT 54.0000 138.3000 54.8000 138.4000 ;
	    RECT 4.4000 137.7000 54.8000 138.3000 ;
	    RECT 4.4000 137.6000 5.2000 137.7000 ;
	    RECT 20.4000 137.6000 21.2000 137.7000 ;
	    RECT 54.0000 137.6000 54.8000 137.7000 ;
	    RECT 58.8000 136.3000 59.6000 136.4000 ;
	    RECT 74.8000 136.3000 75.6000 136.4000 ;
	    RECT 58.8000 135.7000 75.6000 136.3000 ;
	    RECT 58.8000 135.6000 59.6000 135.7000 ;
	    RECT 74.8000 135.6000 75.6000 135.7000 ;
	    RECT 39.6000 134.3000 40.4000 134.4000 ;
	    RECT 49.2000 134.3000 50.0000 134.4000 ;
	    RECT 39.6000 133.7000 50.0000 134.3000 ;
	    RECT 39.6000 133.6000 40.4000 133.7000 ;
	    RECT 49.2000 133.6000 50.0000 133.7000 ;
	    RECT 74.8000 134.3000 75.6000 134.4000 ;
	    RECT 79.6000 134.3000 80.4000 134.4000 ;
	    RECT 74.8000 133.7000 80.4000 134.3000 ;
	    RECT 74.8000 133.6000 75.6000 133.7000 ;
	    RECT 79.6000 133.6000 80.4000 133.7000 ;
	    RECT 81.2000 133.6000 82.0000 134.4000 ;
	    RECT 150.0000 134.3000 150.8000 134.4000 ;
	    RECT 164.4000 134.3000 165.2000 134.4000 ;
	    RECT 150.0000 133.7000 165.2000 134.3000 ;
	    RECT 150.0000 133.6000 150.8000 133.7000 ;
	    RECT 164.4000 133.6000 165.2000 133.7000 ;
	    RECT 17.2000 131.6000 18.0000 132.4000 ;
	    RECT 52.4000 132.3000 53.2000 132.4000 ;
	    RECT 55.6000 132.3000 56.4000 132.4000 ;
	    RECT 60.4000 132.3000 61.2000 132.4000 ;
	    RECT 52.4000 131.7000 61.2000 132.3000 ;
	    RECT 52.4000 131.6000 53.2000 131.7000 ;
	    RECT 55.6000 131.6000 56.4000 131.7000 ;
	    RECT 60.4000 131.6000 61.2000 131.7000 ;
	    RECT 78.0000 132.3000 78.8000 132.4000 ;
	    RECT 82.8000 132.3000 83.6000 132.4000 ;
	    RECT 78.0000 131.7000 83.6000 132.3000 ;
	    RECT 78.0000 131.6000 78.8000 131.7000 ;
	    RECT 82.8000 131.6000 83.6000 131.7000 ;
	    RECT 100.4000 132.3000 101.2000 132.4000 ;
	    RECT 111.6000 132.3000 112.4000 132.4000 ;
	    RECT 100.4000 131.7000 112.4000 132.3000 ;
	    RECT 100.4000 131.6000 101.2000 131.7000 ;
	    RECT 111.6000 131.6000 112.4000 131.7000 ;
	    RECT 158.0000 132.3000 158.8000 132.4000 ;
	    RECT 190.0000 132.3000 190.8000 132.4000 ;
	    RECT 158.0000 131.7000 190.8000 132.3000 ;
	    RECT 158.0000 131.6000 158.8000 131.7000 ;
	    RECT 190.0000 131.6000 190.8000 131.7000 ;
	    RECT 28.4000 128.3000 29.2000 128.4000 ;
	    RECT 39.6000 128.3000 40.4000 128.4000 ;
	    RECT 58.8000 128.3000 59.6000 128.4000 ;
	    RECT 87.6000 128.3000 88.4000 128.4000 ;
	    RECT 28.4000 127.7000 88.4000 128.3000 ;
	    RECT 28.4000 127.6000 29.2000 127.7000 ;
	    RECT 39.6000 127.6000 40.4000 127.7000 ;
	    RECT 58.8000 127.6000 59.6000 127.7000 ;
	    RECT 87.6000 127.6000 88.4000 127.7000 ;
	    RECT 36.4000 124.3000 37.2000 124.4000 ;
	    RECT 54.0000 124.3000 54.8000 124.4000 ;
	    RECT 36.4000 123.7000 54.8000 124.3000 ;
	    RECT 36.4000 123.6000 37.2000 123.7000 ;
	    RECT 54.0000 123.6000 54.8000 123.7000 ;
	    RECT 121.2000 124.3000 122.0000 124.4000 ;
	    RECT 126.0000 124.3000 126.8000 124.4000 ;
	    RECT 143.6000 124.3000 144.4000 124.4000 ;
	    RECT 121.2000 123.7000 144.4000 124.3000 ;
	    RECT 121.2000 123.6000 122.0000 123.7000 ;
	    RECT 126.0000 123.6000 126.8000 123.7000 ;
	    RECT 143.6000 123.6000 144.4000 123.7000 ;
	    RECT 12.4000 122.3000 13.2000 122.4000 ;
	    RECT 15.6000 122.3000 16.4000 122.4000 ;
	    RECT 31.6000 122.3000 32.4000 122.4000 ;
	    RECT 12.4000 121.7000 32.4000 122.3000 ;
	    RECT 12.4000 121.6000 13.2000 121.7000 ;
	    RECT 15.6000 121.6000 16.4000 121.7000 ;
	    RECT 31.6000 121.6000 32.4000 121.7000 ;
	    RECT 194.8000 122.3000 195.6000 122.4000 ;
	    RECT 199.6000 122.3000 200.4000 122.4000 ;
	    RECT 194.8000 121.7000 200.4000 122.3000 ;
	    RECT 194.8000 121.6000 195.6000 121.7000 ;
	    RECT 199.6000 121.6000 200.4000 121.7000 ;
	    RECT 124.4000 118.3000 125.2000 118.4000 ;
	    RECT 143.6000 118.3000 144.4000 118.4000 ;
	    RECT 164.4000 118.3000 165.2000 118.4000 ;
	    RECT 124.4000 117.7000 165.2000 118.3000 ;
	    RECT 124.4000 117.6000 125.2000 117.7000 ;
	    RECT 143.6000 117.6000 144.4000 117.7000 ;
	    RECT 164.4000 117.6000 165.2000 117.7000 ;
	    RECT 130.8000 116.3000 131.6000 116.4000 ;
	    RECT 146.8000 116.3000 147.6000 116.4000 ;
	    RECT 180.4000 116.3000 181.2000 116.4000 ;
	    RECT 183.6000 116.3000 184.4000 116.4000 ;
	    RECT 130.8000 115.7000 184.4000 116.3000 ;
	    RECT 130.8000 115.6000 131.6000 115.7000 ;
	    RECT 146.8000 115.6000 147.6000 115.7000 ;
	    RECT 180.4000 115.6000 181.2000 115.7000 ;
	    RECT 183.6000 115.6000 184.4000 115.7000 ;
	    RECT 79.6000 114.3000 80.4000 114.4000 ;
	    RECT 132.4000 114.3000 133.2000 114.4000 ;
	    RECT 148.4000 114.3000 149.2000 114.4000 ;
	    RECT 79.6000 113.7000 149.2000 114.3000 ;
	    RECT 79.6000 113.6000 80.4000 113.7000 ;
	    RECT 132.4000 113.6000 133.2000 113.7000 ;
	    RECT 148.4000 113.6000 149.2000 113.7000 ;
	    RECT 150.0000 114.3000 150.8000 114.4000 ;
	    RECT 191.6000 114.3000 192.4000 114.4000 ;
	    RECT 150.0000 113.7000 192.4000 114.3000 ;
	    RECT 150.0000 113.6000 150.8000 113.7000 ;
	    RECT 191.6000 113.6000 192.4000 113.7000 ;
	    RECT 17.2000 112.3000 18.0000 112.4000 ;
	    RECT 25.2000 112.3000 26.0000 112.4000 ;
	    RECT 79.7000 112.3000 80.3000 113.6000 ;
	    RECT 17.2000 111.7000 80.3000 112.3000 ;
	    RECT 140.4000 112.3000 141.2000 112.4000 ;
	    RECT 145.2000 112.3000 146.0000 112.4000 ;
	    RECT 174.0000 112.3000 174.8000 112.4000 ;
	    RECT 186.8000 112.3000 187.6000 112.4000 ;
	    RECT 140.4000 111.7000 144.3000 112.3000 ;
	    RECT 17.2000 111.6000 18.0000 111.7000 ;
	    RECT 25.2000 111.6000 26.0000 111.7000 ;
	    RECT 140.4000 111.6000 141.2000 111.7000 ;
	    RECT 36.4000 110.3000 37.2000 110.4000 ;
	    RECT 57.2000 110.3000 58.0000 110.4000 ;
	    RECT 36.4000 109.7000 58.0000 110.3000 ;
	    RECT 36.4000 109.6000 37.2000 109.7000 ;
	    RECT 57.2000 109.6000 58.0000 109.7000 ;
	    RECT 66.8000 110.3000 67.6000 110.4000 ;
	    RECT 98.8000 110.3000 99.6000 110.4000 ;
	    RECT 66.8000 109.7000 99.6000 110.3000 ;
	    RECT 66.8000 109.6000 67.6000 109.7000 ;
	    RECT 98.8000 109.6000 99.6000 109.7000 ;
	    RECT 127.6000 110.3000 128.4000 110.4000 ;
	    RECT 138.8000 110.3000 139.6000 110.4000 ;
	    RECT 142.0000 110.3000 142.8000 110.4000 ;
	    RECT 127.6000 109.7000 142.8000 110.3000 ;
	    RECT 143.7000 110.3000 144.3000 111.7000 ;
	    RECT 145.2000 111.7000 187.6000 112.3000 ;
	    RECT 145.2000 111.6000 146.0000 111.7000 ;
	    RECT 174.0000 111.6000 174.8000 111.7000 ;
	    RECT 186.8000 111.6000 187.6000 111.7000 ;
	    RECT 150.0000 110.3000 150.8000 110.4000 ;
	    RECT 143.7000 109.7000 150.8000 110.3000 ;
	    RECT 127.6000 109.6000 128.4000 109.7000 ;
	    RECT 138.8000 109.6000 139.6000 109.7000 ;
	    RECT 142.0000 109.6000 142.8000 109.7000 ;
	    RECT 150.0000 109.6000 150.8000 109.7000 ;
	    RECT 156.4000 110.3000 157.2000 110.4000 ;
	    RECT 170.8000 110.3000 171.6000 110.4000 ;
	    RECT 156.4000 109.7000 171.6000 110.3000 ;
	    RECT 156.4000 109.6000 157.2000 109.7000 ;
	    RECT 170.8000 109.6000 171.6000 109.7000 ;
	    RECT 182.0000 110.3000 182.8000 110.4000 ;
	    RECT 185.2000 110.3000 186.0000 110.4000 ;
	    RECT 198.0000 110.3000 198.8000 110.4000 ;
	    RECT 182.0000 109.7000 198.8000 110.3000 ;
	    RECT 182.0000 109.6000 182.8000 109.7000 ;
	    RECT 185.2000 109.6000 186.0000 109.7000 ;
	    RECT 198.0000 109.6000 198.8000 109.7000 ;
	    RECT 209.2000 110.3000 210.0000 110.4000 ;
	    RECT 222.0000 110.3000 222.8000 110.4000 ;
	    RECT 209.2000 109.7000 222.8000 110.3000 ;
	    RECT 209.2000 109.6000 210.0000 109.7000 ;
	    RECT 222.0000 109.6000 222.8000 109.7000 ;
	    RECT 10.8000 108.3000 11.6000 108.4000 ;
	    RECT 22.0000 108.3000 22.8000 108.4000 ;
	    RECT 38.0000 108.3000 38.8000 108.4000 ;
	    RECT 169.2000 108.3000 170.0000 108.4000 ;
	    RECT 218.8000 108.3000 219.6000 108.4000 ;
	    RECT 10.8000 107.7000 38.8000 108.3000 ;
	    RECT 10.8000 107.6000 11.6000 107.7000 ;
	    RECT 22.0000 107.6000 22.8000 107.7000 ;
	    RECT 38.0000 107.6000 38.8000 107.7000 ;
	    RECT 153.3000 107.7000 219.6000 108.3000 ;
	    RECT 153.3000 106.4000 153.9000 107.7000 ;
	    RECT 169.2000 107.6000 170.0000 107.7000 ;
	    RECT 218.8000 107.6000 219.6000 107.7000 ;
	    RECT 4.4000 106.3000 5.2000 106.4000 ;
	    RECT 14.0000 106.3000 14.8000 106.4000 ;
	    RECT 4.4000 105.7000 14.8000 106.3000 ;
	    RECT 4.4000 105.6000 5.2000 105.7000 ;
	    RECT 14.0000 105.6000 14.8000 105.7000 ;
	    RECT 22.0000 106.3000 22.8000 106.4000 ;
	    RECT 26.8000 106.3000 27.6000 106.4000 ;
	    RECT 22.0000 105.7000 27.6000 106.3000 ;
	    RECT 22.0000 105.6000 22.8000 105.7000 ;
	    RECT 26.8000 105.6000 27.6000 105.7000 ;
	    RECT 30.0000 106.3000 30.8000 106.4000 ;
	    RECT 44.4000 106.3000 45.2000 106.4000 ;
	    RECT 30.0000 105.7000 45.2000 106.3000 ;
	    RECT 30.0000 105.6000 30.8000 105.7000 ;
	    RECT 44.4000 105.6000 45.2000 105.7000 ;
	    RECT 54.0000 106.3000 54.8000 106.4000 ;
	    RECT 76.4000 106.3000 77.2000 106.4000 ;
	    RECT 79.6000 106.3000 80.4000 106.4000 ;
	    RECT 54.0000 105.7000 80.4000 106.3000 ;
	    RECT 54.0000 105.6000 54.8000 105.7000 ;
	    RECT 76.4000 105.6000 77.2000 105.7000 ;
	    RECT 79.6000 105.6000 80.4000 105.7000 ;
	    RECT 132.4000 106.3000 133.2000 106.4000 ;
	    RECT 153.2000 106.3000 154.0000 106.4000 ;
	    RECT 132.4000 105.7000 154.0000 106.3000 ;
	    RECT 132.4000 105.6000 133.2000 105.7000 ;
	    RECT 153.2000 105.6000 154.0000 105.7000 ;
	    RECT 167.6000 106.3000 168.4000 106.4000 ;
	    RECT 185.2000 106.3000 186.0000 106.4000 ;
	    RECT 167.6000 105.7000 186.0000 106.3000 ;
	    RECT 167.6000 105.6000 168.4000 105.7000 ;
	    RECT 185.2000 105.6000 186.0000 105.7000 ;
	    RECT 204.4000 106.3000 205.2000 106.4000 ;
	    RECT 210.8000 106.3000 211.6000 106.4000 ;
	    RECT 218.8000 106.3000 219.6000 106.4000 ;
	    RECT 204.4000 105.7000 219.6000 106.3000 ;
	    RECT 204.4000 105.6000 205.2000 105.7000 ;
	    RECT 210.8000 105.6000 211.6000 105.7000 ;
	    RECT 218.8000 105.6000 219.6000 105.7000 ;
	    RECT 34.8000 104.3000 35.6000 104.4000 ;
	    RECT 41.2000 104.3000 42.0000 104.4000 ;
	    RECT 34.8000 103.7000 42.0000 104.3000 ;
	    RECT 34.8000 103.6000 35.6000 103.7000 ;
	    RECT 41.2000 103.6000 42.0000 103.7000 ;
	    RECT 135.6000 104.3000 136.4000 104.4000 ;
	    RECT 156.4000 104.3000 157.2000 104.4000 ;
	    RECT 135.6000 103.7000 157.2000 104.3000 ;
	    RECT 135.6000 103.6000 136.4000 103.7000 ;
	    RECT 156.4000 103.6000 157.2000 103.7000 ;
	    RECT 166.0000 104.3000 166.8000 104.4000 ;
	    RECT 175.6000 104.3000 176.4000 104.4000 ;
	    RECT 166.0000 103.7000 176.4000 104.3000 ;
	    RECT 166.0000 103.6000 166.8000 103.7000 ;
	    RECT 175.6000 103.6000 176.4000 103.7000 ;
	    RECT 196.4000 104.3000 197.2000 104.4000 ;
	    RECT 212.4000 104.3000 213.2000 104.4000 ;
	    RECT 196.4000 103.7000 213.2000 104.3000 ;
	    RECT 196.4000 103.6000 197.2000 103.7000 ;
	    RECT 212.4000 103.6000 213.2000 103.7000 ;
	    RECT 78.0000 102.3000 78.8000 102.4000 ;
	    RECT 90.8000 102.3000 91.6000 102.4000 ;
	    RECT 78.0000 101.7000 91.6000 102.3000 ;
	    RECT 78.0000 101.6000 78.8000 101.7000 ;
	    RECT 90.8000 101.6000 91.6000 101.7000 ;
	    RECT 180.4000 102.3000 181.2000 102.4000 ;
	    RECT 209.2000 102.3000 210.0000 102.4000 ;
	    RECT 180.4000 101.7000 210.0000 102.3000 ;
	    RECT 180.4000 101.6000 181.2000 101.7000 ;
	    RECT 209.2000 101.6000 210.0000 101.7000 ;
	    RECT 135.6000 100.3000 136.4000 100.4000 ;
	    RECT 145.2000 100.3000 146.0000 100.4000 ;
	    RECT 135.6000 99.7000 146.0000 100.3000 ;
	    RECT 135.6000 99.6000 136.4000 99.7000 ;
	    RECT 145.2000 99.6000 146.0000 99.7000 ;
	    RECT 38.0000 98.3000 38.8000 98.4000 ;
	    RECT 47.6000 98.3000 48.4000 98.4000 ;
	    RECT 38.0000 97.7000 48.4000 98.3000 ;
	    RECT 38.0000 97.6000 38.8000 97.7000 ;
	    RECT 47.6000 97.6000 48.4000 97.7000 ;
	    RECT 98.8000 98.3000 99.6000 98.4000 ;
	    RECT 108.4000 98.3000 109.2000 98.4000 ;
	    RECT 98.8000 97.7000 109.2000 98.3000 ;
	    RECT 98.8000 97.6000 99.6000 97.7000 ;
	    RECT 108.4000 97.6000 109.2000 97.7000 ;
	    RECT 39.6000 96.3000 40.4000 96.4000 ;
	    RECT 86.0000 96.3000 86.8000 96.4000 ;
	    RECT 110.0000 96.3000 110.8000 96.4000 ;
	    RECT 39.6000 95.7000 46.7000 96.3000 ;
	    RECT 39.6000 95.6000 40.4000 95.7000 ;
	    RECT 46.1000 94.4000 46.7000 95.7000 ;
	    RECT 86.0000 95.7000 110.8000 96.3000 ;
	    RECT 86.0000 95.6000 86.8000 95.7000 ;
	    RECT 110.0000 95.6000 110.8000 95.7000 ;
	    RECT 151.6000 96.3000 152.4000 96.4000 ;
	    RECT 190.0000 96.3000 190.8000 96.4000 ;
	    RECT 151.6000 95.7000 190.8000 96.3000 ;
	    RECT 151.6000 95.6000 152.4000 95.7000 ;
	    RECT 190.0000 95.6000 190.8000 95.7000 ;
	    RECT 28.4000 94.3000 29.2000 94.4000 ;
	    RECT 41.2000 94.3000 42.0000 94.4000 ;
	    RECT 28.4000 93.7000 42.0000 94.3000 ;
	    RECT 28.4000 93.6000 29.2000 93.7000 ;
	    RECT 41.2000 93.6000 42.0000 93.7000 ;
	    RECT 46.0000 94.3000 46.8000 94.4000 ;
	    RECT 57.2000 94.3000 58.0000 94.4000 ;
	    RECT 70.0000 94.3000 70.8000 94.4000 ;
	    RECT 46.0000 93.7000 70.8000 94.3000 ;
	    RECT 46.0000 93.6000 46.8000 93.7000 ;
	    RECT 57.2000 93.6000 58.0000 93.7000 ;
	    RECT 70.0000 93.6000 70.8000 93.7000 ;
	    RECT 74.8000 94.3000 75.6000 94.4000 ;
	    RECT 89.2000 94.3000 90.0000 94.4000 ;
	    RECT 74.8000 93.7000 90.0000 94.3000 ;
	    RECT 74.8000 93.6000 75.6000 93.7000 ;
	    RECT 89.2000 93.6000 90.0000 93.7000 ;
	    RECT 106.8000 94.3000 107.6000 94.4000 ;
	    RECT 113.2000 94.3000 114.0000 94.4000 ;
	    RECT 116.4000 94.3000 117.2000 94.4000 ;
	    RECT 106.8000 93.7000 117.2000 94.3000 ;
	    RECT 106.8000 93.6000 107.6000 93.7000 ;
	    RECT 113.2000 93.6000 114.0000 93.7000 ;
	    RECT 116.4000 93.6000 117.2000 93.7000 ;
	    RECT 154.8000 94.3000 155.6000 94.4000 ;
	    RECT 177.2000 94.3000 178.0000 94.4000 ;
	    RECT 154.8000 93.7000 178.0000 94.3000 ;
	    RECT 154.8000 93.6000 155.6000 93.7000 ;
	    RECT 177.2000 93.6000 178.0000 93.7000 ;
	    RECT 218.8000 94.3000 219.6000 94.4000 ;
	    RECT 220.4000 94.3000 221.2000 94.4000 ;
	    RECT 218.8000 93.7000 221.2000 94.3000 ;
	    RECT 218.8000 93.6000 219.6000 93.7000 ;
	    RECT 220.4000 93.6000 221.2000 93.7000 ;
	    RECT 44.4000 92.3000 45.2000 92.4000 ;
	    RECT 46.0000 92.3000 46.8000 92.4000 ;
	    RECT 58.8000 92.3000 59.6000 92.4000 ;
	    RECT 44.4000 91.7000 59.6000 92.3000 ;
	    RECT 44.4000 91.6000 45.2000 91.7000 ;
	    RECT 46.0000 91.6000 46.8000 91.7000 ;
	    RECT 58.8000 91.6000 59.6000 91.7000 ;
	    RECT 121.2000 92.3000 122.0000 92.4000 ;
	    RECT 126.0000 92.3000 126.8000 92.4000 ;
	    RECT 130.8000 92.3000 131.6000 92.4000 ;
	    RECT 138.8000 92.3000 139.6000 92.4000 ;
	    RECT 121.2000 91.7000 139.6000 92.3000 ;
	    RECT 121.2000 91.6000 122.0000 91.7000 ;
	    RECT 126.0000 91.6000 126.8000 91.7000 ;
	    RECT 130.8000 91.6000 131.6000 91.7000 ;
	    RECT 138.8000 91.6000 139.6000 91.7000 ;
	    RECT 161.2000 92.3000 162.0000 92.4000 ;
	    RECT 177.2000 92.3000 178.0000 92.4000 ;
	    RECT 161.2000 91.7000 178.0000 92.3000 ;
	    RECT 161.2000 91.6000 162.0000 91.7000 ;
	    RECT 177.2000 91.6000 178.0000 91.7000 ;
	    RECT 207.6000 92.3000 208.4000 92.4000 ;
	    RECT 215.6000 92.3000 216.4000 92.4000 ;
	    RECT 207.6000 91.7000 216.4000 92.3000 ;
	    RECT 207.6000 91.6000 208.4000 91.7000 ;
	    RECT 215.6000 91.6000 216.4000 91.7000 ;
	    RECT 217.2000 92.3000 218.0000 92.4000 ;
	    RECT 222.0000 92.3000 222.8000 92.4000 ;
	    RECT 217.2000 91.7000 222.8000 92.3000 ;
	    RECT 217.2000 91.6000 218.0000 91.7000 ;
	    RECT 222.0000 91.6000 222.8000 91.7000 ;
	    RECT 116.4000 90.3000 117.2000 90.4000 ;
	    RECT 143.6000 90.3000 144.4000 90.4000 ;
	    RECT 116.4000 89.7000 144.4000 90.3000 ;
	    RECT 116.4000 89.6000 117.2000 89.7000 ;
	    RECT 143.6000 89.6000 144.4000 89.7000 ;
	    RECT 209.2000 90.3000 210.0000 90.4000 ;
	    RECT 215.6000 90.3000 216.4000 90.4000 ;
	    RECT 209.2000 89.7000 216.4000 90.3000 ;
	    RECT 209.2000 89.6000 210.0000 89.7000 ;
	    RECT 215.6000 89.6000 216.4000 89.7000 ;
	    RECT 202.8000 88.3000 203.6000 88.4000 ;
	    RECT 212.4000 88.3000 213.2000 88.4000 ;
	    RECT 222.0000 88.3000 222.8000 88.4000 ;
	    RECT 202.8000 87.7000 222.8000 88.3000 ;
	    RECT 202.8000 87.6000 203.6000 87.7000 ;
	    RECT 212.4000 87.6000 213.2000 87.7000 ;
	    RECT 222.0000 87.6000 222.8000 87.7000 ;
	    RECT 186.8000 84.3000 187.6000 84.4000 ;
	    RECT 191.6000 84.3000 192.4000 84.4000 ;
	    RECT 186.8000 83.7000 192.4000 84.3000 ;
	    RECT 186.8000 83.6000 187.6000 83.7000 ;
	    RECT 191.6000 83.6000 192.4000 83.7000 ;
	    RECT 103.6000 82.3000 104.4000 82.4000 ;
	    RECT 118.0000 82.3000 118.8000 82.4000 ;
	    RECT 103.6000 81.7000 118.8000 82.3000 ;
	    RECT 103.6000 81.6000 104.4000 81.7000 ;
	    RECT 118.0000 81.6000 118.8000 81.7000 ;
	    RECT 217.2000 82.3000 218.0000 82.4000 ;
	    RECT 223.6000 82.3000 224.4000 82.4000 ;
	    RECT 217.2000 81.7000 224.4000 82.3000 ;
	    RECT 217.2000 81.6000 218.0000 81.7000 ;
	    RECT 223.6000 81.6000 224.4000 81.7000 ;
	    RECT 108.4000 80.3000 109.2000 80.4000 ;
	    RECT 118.0000 80.3000 118.8000 80.4000 ;
	    RECT 108.4000 79.7000 118.8000 80.3000 ;
	    RECT 108.4000 79.6000 109.2000 79.7000 ;
	    RECT 118.0000 79.6000 118.8000 79.7000 ;
	    RECT 206.0000 79.6000 206.8000 80.4000 ;
	    RECT 188.4000 76.3000 189.2000 76.4000 ;
	    RECT 210.8000 76.3000 211.6000 76.4000 ;
	    RECT 188.4000 75.7000 211.6000 76.3000 ;
	    RECT 188.4000 75.6000 189.2000 75.7000 ;
	    RECT 210.8000 75.6000 211.6000 75.7000 ;
	    RECT 42.8000 74.3000 43.6000 74.4000 ;
	    RECT 74.8000 74.3000 75.6000 74.4000 ;
	    RECT 42.8000 73.7000 75.6000 74.3000 ;
	    RECT 42.8000 73.6000 43.6000 73.7000 ;
	    RECT 74.8000 73.6000 75.6000 73.7000 ;
	    RECT 194.8000 74.3000 195.6000 74.4000 ;
	    RECT 206.0000 74.3000 206.8000 74.4000 ;
	    RECT 194.8000 73.7000 206.8000 74.3000 ;
	    RECT 194.8000 73.6000 195.6000 73.7000 ;
	    RECT 206.0000 73.6000 206.8000 73.7000 ;
	    RECT 212.4000 74.3000 213.2000 74.4000 ;
	    RECT 217.2000 74.3000 218.0000 74.4000 ;
	    RECT 212.4000 73.7000 218.0000 74.3000 ;
	    RECT 212.4000 73.6000 213.2000 73.7000 ;
	    RECT 217.2000 73.6000 218.0000 73.7000 ;
	    RECT 54.0000 72.3000 54.8000 72.4000 ;
	    RECT 70.0000 72.3000 70.8000 72.4000 ;
	    RECT 54.0000 71.7000 70.8000 72.3000 ;
	    RECT 54.0000 71.6000 54.8000 71.7000 ;
	    RECT 70.0000 71.6000 70.8000 71.7000 ;
	    RECT 164.4000 72.3000 165.2000 72.4000 ;
	    RECT 185.2000 72.3000 186.0000 72.4000 ;
	    RECT 164.4000 71.7000 186.0000 72.3000 ;
	    RECT 164.4000 71.6000 165.2000 71.7000 ;
	    RECT 185.2000 71.6000 186.0000 71.7000 ;
	    RECT 190.0000 72.3000 190.8000 72.4000 ;
	    RECT 198.0000 72.3000 198.8000 72.4000 ;
	    RECT 209.2000 72.3000 210.0000 72.4000 ;
	    RECT 190.0000 71.7000 210.0000 72.3000 ;
	    RECT 190.0000 71.6000 190.8000 71.7000 ;
	    RECT 198.0000 71.6000 198.8000 71.7000 ;
	    RECT 209.2000 71.6000 210.0000 71.7000 ;
	    RECT 38.0000 70.3000 38.8000 70.4000 ;
	    RECT 46.0000 70.3000 46.8000 70.4000 ;
	    RECT 38.0000 69.7000 46.8000 70.3000 ;
	    RECT 38.0000 69.6000 38.8000 69.7000 ;
	    RECT 46.0000 69.6000 46.8000 69.7000 ;
	    RECT 49.2000 70.3000 50.0000 70.4000 ;
	    RECT 55.6000 70.3000 56.4000 70.4000 ;
	    RECT 49.2000 69.7000 56.4000 70.3000 ;
	    RECT 49.2000 69.6000 50.0000 69.7000 ;
	    RECT 55.6000 69.6000 56.4000 69.7000 ;
	    RECT 78.0000 70.3000 78.8000 70.4000 ;
	    RECT 113.2000 70.3000 114.0000 70.4000 ;
	    RECT 78.0000 69.7000 114.0000 70.3000 ;
	    RECT 78.0000 69.6000 78.8000 69.7000 ;
	    RECT 113.2000 69.6000 114.0000 69.7000 ;
	    RECT 175.6000 70.3000 176.4000 70.4000 ;
	    RECT 185.2000 70.3000 186.0000 70.4000 ;
	    RECT 175.6000 69.7000 186.0000 70.3000 ;
	    RECT 175.6000 69.6000 176.4000 69.7000 ;
	    RECT 185.2000 69.6000 186.0000 69.7000 ;
	    RECT 198.0000 70.3000 198.8000 70.4000 ;
	    RECT 202.8000 70.3000 203.6000 70.4000 ;
	    RECT 198.0000 69.7000 203.6000 70.3000 ;
	    RECT 198.0000 69.6000 198.8000 69.7000 ;
	    RECT 202.8000 69.6000 203.6000 69.7000 ;
	    RECT 207.6000 70.3000 208.4000 70.4000 ;
	    RECT 210.8000 70.3000 211.6000 70.4000 ;
	    RECT 207.6000 69.7000 211.6000 70.3000 ;
	    RECT 207.6000 69.6000 208.4000 69.7000 ;
	    RECT 210.8000 69.6000 211.6000 69.7000 ;
	    RECT 212.4000 70.3000 213.2000 70.4000 ;
	    RECT 217.2000 70.3000 218.0000 70.4000 ;
	    RECT 212.4000 69.7000 218.0000 70.3000 ;
	    RECT 212.4000 69.6000 213.2000 69.7000 ;
	    RECT 217.2000 69.6000 218.0000 69.7000 ;
	    RECT 2.8000 68.3000 3.6000 68.4000 ;
	    RECT 47.6000 68.3000 48.4000 68.4000 ;
	    RECT 2.8000 67.7000 48.4000 68.3000 ;
	    RECT 2.8000 67.6000 3.6000 67.7000 ;
	    RECT 47.6000 67.6000 48.4000 67.7000 ;
	    RECT 50.8000 68.3000 51.6000 68.4000 ;
	    RECT 57.2000 68.3000 58.0000 68.4000 ;
	    RECT 50.8000 67.7000 58.0000 68.3000 ;
	    RECT 50.8000 67.6000 51.6000 67.7000 ;
	    RECT 57.2000 67.6000 58.0000 67.7000 ;
	    RECT 73.2000 68.3000 74.0000 68.4000 ;
	    RECT 94.0000 68.3000 94.8000 68.4000 ;
	    RECT 73.2000 67.7000 94.8000 68.3000 ;
	    RECT 73.2000 67.6000 74.0000 67.7000 ;
	    RECT 94.0000 67.6000 94.8000 67.7000 ;
	    RECT 121.2000 68.3000 122.0000 68.4000 ;
	    RECT 126.0000 68.3000 126.8000 68.4000 ;
	    RECT 129.2000 68.3000 130.0000 68.4000 ;
	    RECT 121.2000 67.7000 130.0000 68.3000 ;
	    RECT 121.2000 67.6000 122.0000 67.7000 ;
	    RECT 126.0000 67.6000 126.8000 67.7000 ;
	    RECT 129.2000 67.6000 130.0000 67.7000 ;
	    RECT 161.2000 68.3000 162.0000 68.4000 ;
	    RECT 164.4000 68.3000 165.2000 68.4000 ;
	    RECT 161.2000 67.7000 165.2000 68.3000 ;
	    RECT 161.2000 67.6000 162.0000 67.7000 ;
	    RECT 164.4000 67.6000 165.2000 67.7000 ;
	    RECT 183.6000 68.3000 184.4000 68.4000 ;
	    RECT 190.0000 68.3000 190.8000 68.4000 ;
	    RECT 183.6000 67.7000 190.8000 68.3000 ;
	    RECT 183.6000 67.6000 184.4000 67.7000 ;
	    RECT 190.0000 67.6000 190.8000 67.7000 ;
	    RECT 54.0000 66.3000 54.8000 66.4000 ;
	    RECT 58.8000 66.3000 59.6000 66.4000 ;
	    RECT 54.0000 65.7000 59.6000 66.3000 ;
	    RECT 54.0000 65.6000 54.8000 65.7000 ;
	    RECT 58.8000 65.6000 59.6000 65.7000 ;
	    RECT 66.8000 66.3000 67.6000 66.4000 ;
	    RECT 79.6000 66.3000 80.4000 66.4000 ;
	    RECT 66.8000 65.7000 80.4000 66.3000 ;
	    RECT 66.8000 65.6000 67.6000 65.7000 ;
	    RECT 79.6000 65.6000 80.4000 65.7000 ;
	    RECT 180.4000 66.3000 181.2000 66.4000 ;
	    RECT 185.2000 66.3000 186.0000 66.4000 ;
	    RECT 196.4000 66.3000 197.2000 66.4000 ;
	    RECT 180.4000 65.7000 197.2000 66.3000 ;
	    RECT 180.4000 65.6000 181.2000 65.7000 ;
	    RECT 185.2000 65.6000 186.0000 65.7000 ;
	    RECT 196.4000 65.6000 197.2000 65.7000 ;
	    RECT 201.2000 66.3000 202.0000 66.4000 ;
	    RECT 202.8000 66.3000 203.6000 66.4000 ;
	    RECT 206.0000 66.3000 206.8000 66.4000 ;
	    RECT 212.4000 66.3000 213.2000 66.4000 ;
	    RECT 201.2000 65.7000 213.2000 66.3000 ;
	    RECT 201.2000 65.6000 202.0000 65.7000 ;
	    RECT 202.8000 65.6000 203.6000 65.7000 ;
	    RECT 206.0000 65.6000 206.8000 65.7000 ;
	    RECT 212.4000 65.6000 213.2000 65.7000 ;
	    RECT 46.0000 64.3000 46.8000 64.4000 ;
	    RECT 55.6000 64.3000 56.4000 64.4000 ;
	    RECT 46.0000 63.7000 56.4000 64.3000 ;
	    RECT 46.0000 63.6000 46.8000 63.7000 ;
	    RECT 55.6000 63.6000 56.4000 63.7000 ;
	    RECT 74.8000 64.3000 75.6000 64.4000 ;
	    RECT 97.2000 64.3000 98.0000 64.4000 ;
	    RECT 74.8000 63.7000 98.0000 64.3000 ;
	    RECT 74.8000 63.6000 75.6000 63.7000 ;
	    RECT 97.2000 63.6000 98.0000 63.7000 ;
	    RECT 142.0000 64.3000 142.8000 64.4000 ;
	    RECT 153.2000 64.3000 154.0000 64.4000 ;
	    RECT 164.4000 64.3000 165.2000 64.4000 ;
	    RECT 142.0000 63.7000 165.2000 64.3000 ;
	    RECT 142.0000 63.6000 142.8000 63.7000 ;
	    RECT 153.2000 63.6000 154.0000 63.7000 ;
	    RECT 164.4000 63.6000 165.2000 63.7000 ;
	    RECT 180.4000 64.3000 181.2000 64.4000 ;
	    RECT 186.8000 64.3000 187.6000 64.4000 ;
	    RECT 180.4000 63.7000 187.6000 64.3000 ;
	    RECT 180.4000 63.6000 181.2000 63.7000 ;
	    RECT 186.8000 63.6000 187.6000 63.7000 ;
	    RECT 215.6000 64.3000 216.4000 64.4000 ;
	    RECT 218.8000 64.3000 219.6000 64.4000 ;
	    RECT 215.6000 63.7000 219.6000 64.3000 ;
	    RECT 215.6000 63.6000 216.4000 63.7000 ;
	    RECT 218.8000 63.6000 219.6000 63.7000 ;
	    RECT 22.0000 62.3000 22.8000 62.4000 ;
	    RECT 26.8000 62.3000 27.6000 62.4000 ;
	    RECT 22.0000 61.7000 27.6000 62.3000 ;
	    RECT 22.0000 61.6000 22.8000 61.7000 ;
	    RECT 26.8000 61.6000 27.6000 61.7000 ;
	    RECT 28.4000 62.3000 29.2000 62.4000 ;
	    RECT 42.8000 62.3000 43.6000 62.4000 ;
	    RECT 28.4000 61.7000 43.6000 62.3000 ;
	    RECT 28.4000 61.6000 29.2000 61.7000 ;
	    RECT 42.8000 61.6000 43.6000 61.7000 ;
	    RECT 103.6000 62.3000 104.4000 62.4000 ;
	    RECT 124.4000 62.3000 125.2000 62.4000 ;
	    RECT 103.6000 61.7000 125.2000 62.3000 ;
	    RECT 103.6000 61.6000 104.4000 61.7000 ;
	    RECT 124.4000 61.6000 125.2000 61.7000 ;
	    RECT 22.0000 60.3000 22.8000 60.4000 ;
	    RECT 36.4000 60.3000 37.2000 60.4000 ;
	    RECT 22.0000 59.7000 37.2000 60.3000 ;
	    RECT 22.0000 59.6000 22.8000 59.7000 ;
	    RECT 36.4000 59.6000 37.2000 59.7000 ;
	    RECT 18.8000 58.3000 19.6000 58.4000 ;
	    RECT 23.6000 58.3000 24.4000 58.4000 ;
	    RECT 18.8000 57.7000 24.4000 58.3000 ;
	    RECT 18.8000 57.6000 19.6000 57.7000 ;
	    RECT 23.6000 57.6000 24.4000 57.7000 ;
	    RECT 34.8000 58.3000 35.6000 58.4000 ;
	    RECT 41.2000 58.3000 42.0000 58.4000 ;
	    RECT 34.8000 57.7000 42.0000 58.3000 ;
	    RECT 34.8000 57.6000 35.6000 57.7000 ;
	    RECT 41.2000 57.6000 42.0000 57.7000 ;
	    RECT 164.4000 58.3000 165.2000 58.4000 ;
	    RECT 190.0000 58.3000 190.8000 58.4000 ;
	    RECT 199.6000 58.3000 200.4000 58.4000 ;
	    RECT 164.4000 57.7000 200.4000 58.3000 ;
	    RECT 164.4000 57.6000 165.2000 57.7000 ;
	    RECT 190.0000 57.6000 190.8000 57.7000 ;
	    RECT 199.6000 57.6000 200.4000 57.7000 ;
	    RECT 4.4000 56.3000 5.2000 56.4000 ;
	    RECT 22.0000 56.3000 22.8000 56.4000 ;
	    RECT 4.4000 55.7000 22.8000 56.3000 ;
	    RECT 4.4000 55.6000 5.2000 55.7000 ;
	    RECT 22.0000 55.6000 22.8000 55.7000 ;
	    RECT 31.6000 56.3000 32.4000 56.4000 ;
	    RECT 36.4000 56.3000 37.2000 56.4000 ;
	    RECT 52.4000 56.3000 53.2000 56.4000 ;
	    RECT 31.6000 55.7000 53.2000 56.3000 ;
	    RECT 31.6000 55.6000 32.4000 55.7000 ;
	    RECT 36.4000 55.6000 37.2000 55.7000 ;
	    RECT 52.4000 55.6000 53.2000 55.7000 ;
	    RECT 102.0000 56.3000 102.8000 56.4000 ;
	    RECT 103.6000 56.3000 104.4000 56.4000 ;
	    RECT 102.0000 55.7000 104.4000 56.3000 ;
	    RECT 102.0000 55.6000 102.8000 55.7000 ;
	    RECT 103.6000 55.6000 104.4000 55.7000 ;
	    RECT 210.8000 56.3000 211.6000 56.4000 ;
	    RECT 217.2000 56.3000 218.0000 56.4000 ;
	    RECT 210.8000 55.7000 218.0000 56.3000 ;
	    RECT 210.8000 55.6000 211.6000 55.7000 ;
	    RECT 217.2000 55.6000 218.0000 55.7000 ;
	    RECT 9.2000 54.3000 10.0000 54.4000 ;
	    RECT 38.0000 54.3000 38.8000 54.4000 ;
	    RECT 9.2000 53.7000 38.8000 54.3000 ;
	    RECT 9.2000 53.6000 10.0000 53.7000 ;
	    RECT 38.0000 53.6000 38.8000 53.7000 ;
	    RECT 100.4000 54.3000 101.2000 54.4000 ;
	    RECT 110.0000 54.3000 110.8000 54.4000 ;
	    RECT 142.0000 54.3000 142.8000 54.4000 ;
	    RECT 100.4000 53.7000 142.8000 54.3000 ;
	    RECT 100.4000 53.6000 101.2000 53.7000 ;
	    RECT 110.0000 53.6000 110.8000 53.7000 ;
	    RECT 142.0000 53.6000 142.8000 53.7000 ;
	    RECT 145.2000 54.3000 146.0000 54.4000 ;
	    RECT 167.6000 54.3000 168.4000 54.4000 ;
	    RECT 145.2000 53.7000 168.4000 54.3000 ;
	    RECT 145.2000 53.6000 146.0000 53.7000 ;
	    RECT 167.6000 53.6000 168.4000 53.7000 ;
	    RECT 170.8000 54.3000 171.6000 54.4000 ;
	    RECT 177.2000 54.3000 178.0000 54.4000 ;
	    RECT 170.8000 53.7000 178.0000 54.3000 ;
	    RECT 170.8000 53.6000 171.6000 53.7000 ;
	    RECT 177.2000 53.6000 178.0000 53.7000 ;
	    RECT 183.6000 54.3000 184.4000 54.4000 ;
	    RECT 198.0000 54.3000 198.8000 54.4000 ;
	    RECT 183.6000 53.7000 198.8000 54.3000 ;
	    RECT 183.6000 53.6000 184.4000 53.7000 ;
	    RECT 198.0000 53.6000 198.8000 53.7000 ;
	    RECT 204.4000 54.3000 205.2000 54.4000 ;
	    RECT 214.0000 54.3000 214.8000 54.4000 ;
	    RECT 204.4000 53.7000 214.8000 54.3000 ;
	    RECT 204.4000 53.6000 205.2000 53.7000 ;
	    RECT 214.0000 53.6000 214.8000 53.7000 ;
	    RECT 2.8000 52.3000 3.6000 52.4000 ;
	    RECT 12.4000 52.3000 13.2000 52.4000 ;
	    RECT 2.8000 51.7000 13.2000 52.3000 ;
	    RECT 2.8000 51.6000 3.6000 51.7000 ;
	    RECT 12.4000 51.6000 13.2000 51.7000 ;
	    RECT 17.2000 52.3000 18.0000 52.4000 ;
	    RECT 18.8000 52.3000 19.6000 52.4000 ;
	    RECT 50.8000 52.3000 51.6000 52.4000 ;
	    RECT 17.2000 51.7000 51.6000 52.3000 ;
	    RECT 17.2000 51.6000 18.0000 51.7000 ;
	    RECT 18.8000 51.6000 19.6000 51.7000 ;
	    RECT 50.8000 51.6000 51.6000 51.7000 ;
	    RECT 57.2000 52.3000 58.0000 52.4000 ;
	    RECT 70.0000 52.3000 70.8000 52.4000 ;
	    RECT 57.2000 51.7000 70.8000 52.3000 ;
	    RECT 57.2000 51.6000 58.0000 51.7000 ;
	    RECT 70.0000 51.6000 70.8000 51.7000 ;
	    RECT 111.6000 52.3000 112.4000 52.4000 ;
	    RECT 121.2000 52.3000 122.0000 52.4000 ;
	    RECT 111.6000 51.7000 122.0000 52.3000 ;
	    RECT 111.6000 51.6000 112.4000 51.7000 ;
	    RECT 121.2000 51.6000 122.0000 51.7000 ;
	    RECT 127.6000 52.3000 128.4000 52.4000 ;
	    RECT 166.0000 52.3000 166.8000 52.4000 ;
	    RECT 127.6000 51.7000 166.8000 52.3000 ;
	    RECT 127.6000 51.6000 128.4000 51.7000 ;
	    RECT 166.0000 51.6000 166.8000 51.7000 ;
	    RECT 177.2000 52.3000 178.0000 52.4000 ;
	    RECT 182.0000 52.3000 182.8000 52.4000 ;
	    RECT 186.8000 52.3000 187.6000 52.4000 ;
	    RECT 177.2000 51.7000 187.6000 52.3000 ;
	    RECT 198.1000 52.3000 198.7000 53.6000 ;
	    RECT 204.4000 52.3000 205.2000 52.4000 ;
	    RECT 206.0000 52.3000 206.8000 52.4000 ;
	    RECT 198.1000 51.7000 206.8000 52.3000 ;
	    RECT 177.2000 51.6000 178.0000 51.7000 ;
	    RECT 182.0000 51.6000 182.8000 51.7000 ;
	    RECT 186.8000 51.6000 187.6000 51.7000 ;
	    RECT 204.4000 51.6000 205.2000 51.7000 ;
	    RECT 206.0000 51.6000 206.8000 51.7000 ;
	    RECT 17.2000 50.3000 18.0000 50.4000 ;
	    RECT 20.4000 50.3000 21.2000 50.4000 ;
	    RECT 17.2000 49.7000 21.2000 50.3000 ;
	    RECT 17.2000 49.6000 18.0000 49.7000 ;
	    RECT 20.4000 49.6000 21.2000 49.7000 ;
	    RECT 106.8000 50.3000 107.6000 50.4000 ;
	    RECT 113.2000 50.3000 114.0000 50.4000 ;
	    RECT 119.6000 50.3000 120.4000 50.4000 ;
	    RECT 106.8000 49.7000 120.4000 50.3000 ;
	    RECT 106.8000 49.6000 107.6000 49.7000 ;
	    RECT 113.2000 49.6000 114.0000 49.7000 ;
	    RECT 119.6000 49.6000 120.4000 49.7000 ;
	    RECT 121.2000 50.3000 122.0000 50.4000 ;
	    RECT 183.6000 50.3000 184.4000 50.4000 ;
	    RECT 121.2000 49.7000 184.4000 50.3000 ;
	    RECT 121.2000 49.6000 122.0000 49.7000 ;
	    RECT 183.6000 49.6000 184.4000 49.7000 ;
	    RECT 23.6000 48.3000 24.4000 48.4000 ;
	    RECT 30.0000 48.3000 30.8000 48.4000 ;
	    RECT 60.4000 48.3000 61.2000 48.4000 ;
	    RECT 90.8000 48.3000 91.6000 48.4000 ;
	    RECT 23.6000 47.7000 91.6000 48.3000 ;
	    RECT 23.6000 47.6000 24.4000 47.7000 ;
	    RECT 30.0000 47.6000 30.8000 47.7000 ;
	    RECT 60.4000 47.6000 61.2000 47.7000 ;
	    RECT 90.8000 47.6000 91.6000 47.7000 ;
	    RECT 114.8000 48.3000 115.6000 48.4000 ;
	    RECT 134.0000 48.3000 134.8000 48.4000 ;
	    RECT 114.8000 47.7000 134.8000 48.3000 ;
	    RECT 114.8000 47.6000 115.6000 47.7000 ;
	    RECT 134.0000 47.6000 134.8000 47.7000 ;
	    RECT 180.4000 48.3000 181.2000 48.4000 ;
	    RECT 188.4000 48.3000 189.2000 48.4000 ;
	    RECT 180.4000 47.7000 189.2000 48.3000 ;
	    RECT 180.4000 47.6000 181.2000 47.7000 ;
	    RECT 188.4000 47.6000 189.2000 47.7000 ;
	    RECT 121.2000 46.3000 122.0000 46.4000 ;
	    RECT 172.4000 46.3000 173.2000 46.4000 ;
	    RECT 121.2000 45.7000 173.2000 46.3000 ;
	    RECT 121.2000 45.6000 122.0000 45.7000 ;
	    RECT 172.4000 45.6000 173.2000 45.7000 ;
	    RECT 169.2000 44.3000 170.0000 44.4000 ;
	    RECT 210.8000 44.3000 211.6000 44.4000 ;
	    RECT 169.2000 43.7000 211.6000 44.3000 ;
	    RECT 169.2000 43.6000 170.0000 43.7000 ;
	    RECT 210.8000 43.6000 211.6000 43.7000 ;
	    RECT 100.4000 42.3000 101.2000 42.4000 ;
	    RECT 122.8000 42.3000 123.6000 42.4000 ;
	    RECT 100.4000 41.7000 123.6000 42.3000 ;
	    RECT 100.4000 41.6000 101.2000 41.7000 ;
	    RECT 122.8000 41.6000 123.6000 41.7000 ;
	    RECT 25.2000 40.3000 26.0000 40.4000 ;
	    RECT 34.8000 40.3000 35.6000 40.4000 ;
	    RECT 25.2000 39.7000 35.6000 40.3000 ;
	    RECT 25.2000 39.6000 26.0000 39.7000 ;
	    RECT 34.8000 39.6000 35.6000 39.7000 ;
	    RECT 6.0000 38.3000 6.8000 38.4000 ;
	    RECT 9.2000 38.3000 10.0000 38.4000 ;
	    RECT 6.0000 37.7000 10.0000 38.3000 ;
	    RECT 6.0000 37.6000 6.8000 37.7000 ;
	    RECT 9.2000 37.6000 10.0000 37.7000 ;
	    RECT 100.4000 36.3000 101.2000 36.4000 ;
	    RECT 84.5000 35.7000 101.2000 36.3000 ;
	    RECT 84.5000 34.4000 85.1000 35.7000 ;
	    RECT 100.4000 35.6000 101.2000 35.7000 ;
	    RECT 105.2000 36.3000 106.0000 36.4000 ;
	    RECT 108.4000 36.3000 109.2000 36.4000 ;
	    RECT 116.4000 36.3000 117.2000 36.4000 ;
	    RECT 105.2000 35.7000 117.2000 36.3000 ;
	    RECT 105.2000 35.6000 106.0000 35.7000 ;
	    RECT 108.4000 35.6000 109.2000 35.7000 ;
	    RECT 116.4000 35.6000 117.2000 35.7000 ;
	    RECT 190.0000 36.3000 190.8000 36.4000 ;
	    RECT 194.8000 36.3000 195.6000 36.4000 ;
	    RECT 190.0000 35.7000 195.6000 36.3000 ;
	    RECT 190.0000 35.6000 190.8000 35.7000 ;
	    RECT 194.8000 35.6000 195.6000 35.7000 ;
	    RECT 55.6000 33.6000 56.4000 34.4000 ;
	    RECT 71.6000 34.3000 72.4000 34.4000 ;
	    RECT 79.6000 34.3000 80.4000 34.4000 ;
	    RECT 84.4000 34.3000 85.2000 34.4000 ;
	    RECT 71.6000 33.7000 85.2000 34.3000 ;
	    RECT 71.6000 33.6000 72.4000 33.7000 ;
	    RECT 79.6000 33.6000 80.4000 33.7000 ;
	    RECT 84.4000 33.6000 85.2000 33.7000 ;
	    RECT 92.4000 34.3000 93.2000 34.4000 ;
	    RECT 113.2000 34.3000 114.0000 34.4000 ;
	    RECT 92.4000 33.7000 114.0000 34.3000 ;
	    RECT 92.4000 33.6000 93.2000 33.7000 ;
	    RECT 113.2000 33.6000 114.0000 33.7000 ;
	    RECT 116.4000 34.3000 117.2000 34.4000 ;
	    RECT 193.2000 34.3000 194.0000 34.4000 ;
	    RECT 116.4000 33.7000 194.0000 34.3000 ;
	    RECT 116.4000 33.6000 117.2000 33.7000 ;
	    RECT 193.2000 33.6000 194.0000 33.7000 ;
	    RECT 194.8000 34.3000 195.6000 34.4000 ;
	    RECT 215.6000 34.3000 216.4000 34.4000 ;
	    RECT 194.8000 33.7000 216.4000 34.3000 ;
	    RECT 194.8000 33.6000 195.6000 33.7000 ;
	    RECT 215.6000 33.6000 216.4000 33.7000 ;
	    RECT 22.0000 32.3000 22.8000 32.4000 ;
	    RECT 23.6000 32.3000 24.4000 32.4000 ;
	    RECT 55.6000 32.3000 56.4000 32.4000 ;
	    RECT 74.8000 32.3000 75.6000 32.4000 ;
	    RECT 22.0000 31.7000 75.6000 32.3000 ;
	    RECT 22.0000 31.6000 22.8000 31.7000 ;
	    RECT 23.6000 31.6000 24.4000 31.7000 ;
	    RECT 55.6000 31.6000 56.4000 31.7000 ;
	    RECT 74.8000 31.6000 75.6000 31.7000 ;
	    RECT 76.4000 32.3000 77.2000 32.4000 ;
	    RECT 79.6000 32.3000 80.4000 32.4000 ;
	    RECT 111.6000 32.3000 112.4000 32.4000 ;
	    RECT 76.4000 31.7000 112.4000 32.3000 ;
	    RECT 76.4000 31.6000 77.2000 31.7000 ;
	    RECT 79.6000 31.6000 80.4000 31.7000 ;
	    RECT 111.6000 31.6000 112.4000 31.7000 ;
	    RECT 191.6000 32.3000 192.4000 32.4000 ;
	    RECT 198.0000 32.3000 198.8000 32.4000 ;
	    RECT 191.6000 31.7000 198.8000 32.3000 ;
	    RECT 191.6000 31.6000 192.4000 31.7000 ;
	    RECT 198.0000 31.6000 198.8000 31.7000 ;
	    RECT 63.6000 30.3000 64.4000 30.4000 ;
	    RECT 82.8000 30.3000 83.6000 30.4000 ;
	    RECT 63.6000 29.7000 83.6000 30.3000 ;
	    RECT 63.6000 29.6000 64.4000 29.7000 ;
	    RECT 82.8000 29.6000 83.6000 29.7000 ;
	    RECT 98.8000 30.3000 99.6000 30.4000 ;
	    RECT 102.0000 30.3000 102.8000 30.4000 ;
	    RECT 98.8000 29.7000 102.8000 30.3000 ;
	    RECT 98.8000 29.6000 99.6000 29.7000 ;
	    RECT 102.0000 29.6000 102.8000 29.7000 ;
	    RECT 201.2000 30.3000 202.0000 30.4000 ;
	    RECT 202.8000 30.3000 203.6000 30.4000 ;
	    RECT 206.0000 30.3000 206.8000 30.4000 ;
	    RECT 201.2000 29.7000 206.8000 30.3000 ;
	    RECT 201.2000 29.6000 202.0000 29.7000 ;
	    RECT 202.8000 29.6000 203.6000 29.7000 ;
	    RECT 206.0000 29.6000 206.8000 29.7000 ;
	    RECT 210.8000 30.3000 211.6000 30.4000 ;
	    RECT 217.2000 30.3000 218.0000 30.4000 ;
	    RECT 210.8000 29.7000 218.0000 30.3000 ;
	    RECT 210.8000 29.6000 211.6000 29.7000 ;
	    RECT 217.2000 29.6000 218.0000 29.7000 ;
	    RECT 52.4000 28.3000 53.2000 28.4000 ;
	    RECT 81.2000 28.3000 82.0000 28.4000 ;
	    RECT 52.4000 27.7000 82.0000 28.3000 ;
	    RECT 52.4000 27.6000 53.2000 27.7000 ;
	    RECT 81.2000 27.6000 82.0000 27.7000 ;
	    RECT 95.6000 28.3000 96.4000 28.4000 ;
	    RECT 110.0000 28.3000 110.8000 28.4000 ;
	    RECT 95.6000 27.7000 110.8000 28.3000 ;
	    RECT 95.6000 27.6000 96.4000 27.7000 ;
	    RECT 110.0000 27.6000 110.8000 27.7000 ;
	    RECT 111.6000 28.3000 112.4000 28.4000 ;
	    RECT 161.2000 28.3000 162.0000 28.4000 ;
	    RECT 111.6000 27.7000 162.0000 28.3000 ;
	    RECT 111.6000 27.6000 112.4000 27.7000 ;
	    RECT 161.2000 27.6000 162.0000 27.7000 ;
	    RECT 167.6000 28.3000 168.4000 28.4000 ;
	    RECT 175.6000 28.3000 176.4000 28.4000 ;
	    RECT 167.6000 27.7000 176.4000 28.3000 ;
	    RECT 167.6000 27.6000 168.4000 27.7000 ;
	    RECT 175.6000 27.6000 176.4000 27.7000 ;
	    RECT 177.2000 28.3000 178.0000 28.4000 ;
	    RECT 180.4000 28.3000 181.2000 28.4000 ;
	    RECT 177.2000 27.7000 181.2000 28.3000 ;
	    RECT 177.2000 27.6000 178.0000 27.7000 ;
	    RECT 180.4000 27.6000 181.2000 27.7000 ;
	    RECT 89.2000 26.3000 90.0000 26.4000 ;
	    RECT 97.2000 26.3000 98.0000 26.4000 ;
	    RECT 89.2000 25.7000 98.0000 26.3000 ;
	    RECT 89.2000 25.6000 90.0000 25.7000 ;
	    RECT 97.2000 25.6000 98.0000 25.7000 ;
	    RECT 110.0000 26.3000 110.8000 26.4000 ;
	    RECT 118.0000 26.3000 118.8000 26.4000 ;
	    RECT 110.0000 25.7000 118.8000 26.3000 ;
	    RECT 110.0000 25.6000 110.8000 25.7000 ;
	    RECT 118.0000 25.6000 118.8000 25.7000 ;
	    RECT 119.6000 26.3000 120.4000 26.4000 ;
	    RECT 162.8000 26.3000 163.6000 26.4000 ;
	    RECT 169.2000 26.3000 170.0000 26.4000 ;
	    RECT 119.6000 25.7000 170.0000 26.3000 ;
	    RECT 119.6000 25.6000 120.4000 25.7000 ;
	    RECT 162.8000 25.6000 163.6000 25.7000 ;
	    RECT 169.2000 25.6000 170.0000 25.7000 ;
	    RECT 170.8000 26.3000 171.6000 26.4000 ;
	    RECT 177.2000 26.3000 178.0000 26.4000 ;
	    RECT 188.4000 26.3000 189.2000 26.4000 ;
	    RECT 170.8000 25.7000 189.2000 26.3000 ;
	    RECT 170.8000 25.6000 171.6000 25.7000 ;
	    RECT 177.2000 25.6000 178.0000 25.7000 ;
	    RECT 188.4000 25.6000 189.2000 25.7000 ;
	    RECT 199.6000 26.3000 200.4000 26.4000 ;
	    RECT 204.4000 26.3000 205.2000 26.4000 ;
	    RECT 199.6000 25.7000 205.2000 26.3000 ;
	    RECT 199.6000 25.6000 200.4000 25.7000 ;
	    RECT 204.4000 25.6000 205.2000 25.7000 ;
	    RECT 142.0000 24.3000 142.8000 24.4000 ;
	    RECT 186.8000 24.3000 187.6000 24.4000 ;
	    RECT 142.0000 23.7000 187.6000 24.3000 ;
	    RECT 142.0000 23.6000 142.8000 23.7000 ;
	    RECT 186.8000 23.6000 187.6000 23.7000 ;
	    RECT 193.2000 24.3000 194.0000 24.4000 ;
	    RECT 209.2000 24.3000 210.0000 24.4000 ;
	    RECT 193.2000 23.7000 210.0000 24.3000 ;
	    RECT 193.2000 23.6000 194.0000 23.7000 ;
	    RECT 209.2000 23.6000 210.0000 23.7000 ;
	    RECT 182.0000 22.3000 182.8000 22.4000 ;
	    RECT 220.4000 22.3000 221.2000 22.4000 ;
	    RECT 182.0000 21.7000 221.2000 22.3000 ;
	    RECT 182.0000 21.6000 182.8000 21.7000 ;
	    RECT 220.4000 21.6000 221.2000 21.7000 ;
	    RECT 161.2000 20.3000 162.0000 20.4000 ;
	    RECT 185.2000 20.3000 186.0000 20.4000 ;
	    RECT 161.2000 19.7000 186.0000 20.3000 ;
	    RECT 161.2000 19.6000 162.0000 19.7000 ;
	    RECT 185.2000 19.6000 186.0000 19.7000 ;
	    RECT 1.2000 18.3000 2.0000 18.4000 ;
	    RECT 7.6000 18.3000 8.4000 18.4000 ;
	    RECT 1.2000 17.7000 8.4000 18.3000 ;
	    RECT 1.2000 17.6000 2.0000 17.7000 ;
	    RECT 7.6000 17.6000 8.4000 17.7000 ;
	    RECT 126.0000 18.3000 126.8000 18.4000 ;
	    RECT 130.8000 18.3000 131.6000 18.4000 ;
	    RECT 135.6000 18.3000 136.4000 18.4000 ;
	    RECT 126.0000 17.7000 136.4000 18.3000 ;
	    RECT 126.0000 17.6000 126.8000 17.7000 ;
	    RECT 130.8000 17.6000 131.6000 17.7000 ;
	    RECT 135.6000 17.6000 136.4000 17.7000 ;
	    RECT 137.2000 18.3000 138.0000 18.4000 ;
	    RECT 146.8000 18.3000 147.6000 18.4000 ;
	    RECT 137.2000 17.7000 147.6000 18.3000 ;
	    RECT 137.2000 17.6000 138.0000 17.7000 ;
	    RECT 146.8000 17.6000 147.6000 17.7000 ;
	    RECT 156.4000 18.3000 157.2000 18.4000 ;
	    RECT 210.8000 18.3000 211.6000 18.4000 ;
	    RECT 156.4000 17.7000 211.6000 18.3000 ;
	    RECT 156.4000 17.6000 157.2000 17.7000 ;
	    RECT 210.8000 17.6000 211.6000 17.7000 ;
	    RECT 126.0000 16.3000 126.8000 16.4000 ;
	    RECT 129.2000 16.3000 130.0000 16.4000 ;
	    RECT 126.0000 15.7000 130.0000 16.3000 ;
	    RECT 126.0000 15.6000 126.8000 15.7000 ;
	    RECT 129.2000 15.6000 130.0000 15.7000 ;
	    RECT 145.2000 16.3000 146.0000 16.4000 ;
	    RECT 153.2000 16.3000 154.0000 16.4000 ;
	    RECT 145.2000 15.7000 154.0000 16.3000 ;
	    RECT 145.2000 15.6000 146.0000 15.7000 ;
	    RECT 153.2000 15.6000 154.0000 15.7000 ;
	    RECT 206.0000 16.3000 206.8000 16.4000 ;
	    RECT 218.8000 16.3000 219.6000 16.4000 ;
	    RECT 206.0000 15.7000 219.6000 16.3000 ;
	    RECT 206.0000 15.6000 206.8000 15.7000 ;
	    RECT 218.8000 15.6000 219.6000 15.7000 ;
	    RECT 14.0000 14.3000 14.8000 14.4000 ;
	    RECT 26.8000 14.3000 27.6000 14.4000 ;
	    RECT 14.0000 13.7000 27.6000 14.3000 ;
	    RECT 14.0000 13.6000 14.8000 13.7000 ;
	    RECT 26.8000 13.6000 27.6000 13.7000 ;
	    RECT 54.0000 14.3000 54.8000 14.4000 ;
	    RECT 55.6000 14.3000 56.4000 14.4000 ;
	    RECT 54.0000 13.7000 56.4000 14.3000 ;
	    RECT 54.0000 13.6000 54.8000 13.7000 ;
	    RECT 55.6000 13.6000 56.4000 13.7000 ;
	    RECT 90.8000 14.3000 91.6000 14.4000 ;
	    RECT 140.4000 14.3000 141.2000 14.4000 ;
	    RECT 90.8000 13.7000 141.2000 14.3000 ;
	    RECT 90.8000 13.6000 91.6000 13.7000 ;
	    RECT 140.4000 13.6000 141.2000 13.7000 ;
	    RECT 146.8000 14.3000 147.6000 14.4000 ;
	    RECT 172.4000 14.3000 173.2000 14.4000 ;
	    RECT 146.8000 13.7000 173.2000 14.3000 ;
	    RECT 146.8000 13.6000 147.6000 13.7000 ;
	    RECT 172.4000 13.6000 173.2000 13.7000 ;
	    RECT 36.4000 12.3000 37.2000 12.4000 ;
	    RECT 44.4000 12.3000 45.2000 12.4000 ;
	    RECT 36.4000 11.7000 45.2000 12.3000 ;
	    RECT 36.4000 11.6000 37.2000 11.7000 ;
	    RECT 44.4000 11.6000 45.2000 11.7000 ;
	    RECT 121.2000 12.3000 122.0000 12.4000 ;
	    RECT 134.0000 12.3000 134.8000 12.4000 ;
	    RECT 121.2000 11.7000 134.8000 12.3000 ;
	    RECT 121.2000 11.6000 122.0000 11.7000 ;
	    RECT 134.0000 11.6000 134.8000 11.7000 ;
	    RECT 135.6000 12.3000 136.4000 12.4000 ;
	    RECT 142.0000 12.3000 142.8000 12.4000 ;
	    RECT 135.6000 11.7000 142.8000 12.3000 ;
	    RECT 135.6000 11.6000 136.4000 11.7000 ;
	    RECT 142.0000 11.6000 142.8000 11.7000 ;
	    RECT 151.6000 12.3000 152.4000 12.4000 ;
	    RECT 178.8000 12.3000 179.6000 12.4000 ;
	    RECT 151.6000 11.7000 179.6000 12.3000 ;
	    RECT 151.6000 11.6000 152.4000 11.7000 ;
	    RECT 178.8000 11.6000 179.6000 11.7000 ;
	    RECT 151.6000 10.3000 152.4000 10.4000 ;
	    RECT 161.2000 10.3000 162.0000 10.4000 ;
	    RECT 151.6000 9.7000 162.0000 10.3000 ;
	    RECT 151.6000 9.6000 152.4000 9.7000 ;
	    RECT 161.2000 9.6000 162.0000 9.7000 ;
	    RECT 209.2000 10.3000 210.0000 10.4000 ;
	    RECT 212.4000 10.3000 213.2000 10.4000 ;
	    RECT 209.2000 9.7000 213.2000 10.3000 ;
	    RECT 209.2000 9.6000 210.0000 9.7000 ;
	    RECT 212.4000 9.6000 213.2000 9.7000 ;
         LAYER metal4 ;
	    RECT 17.0000 51.4000 18.2000 160.6000 ;
	    RECT 39.4000 127.4000 40.6000 148.6000 ;
	    RECT 81.0000 133.4000 82.2000 182.6000 ;
	    RECT 151.4000 181.4000 152.6000 188.6000 ;
	    RECT 116.2000 93.4000 117.4000 170.6000 ;
	    RECT 23.4000 31.4000 24.6000 58.6000 ;
	    RECT 103.4000 55.4000 104.6000 82.6000 ;
	    RECT 164.2000 67.4000 165.4000 72.6000 ;
	    RECT 180.2000 65.4000 181.4000 116.6000 ;
	    RECT 55.4000 13.4000 56.6000 34.6000 ;
	    RECT 202.6000 29.4000 203.8000 88.6000 ;
	    RECT 205.8000 51.4000 207.0000 80.6000 ;
	    RECT 218.6000 63.4000 219.8000 94.6000 ;
   END
END map9v3
