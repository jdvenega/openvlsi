magic
tech scmos
magscale 1 2
timestamp 1560284232
<< metal1 >>
rect 632 2006 638 2014
rect 646 2006 652 2014
rect 660 2006 666 2014
rect 674 2006 680 2014
rect 1604 1977 1619 1983
rect 45 1897 82 1903
rect 445 1897 530 1903
rect 1021 1897 1043 1903
rect 2109 1897 2131 1903
rect 1069 1877 1084 1883
rect 2052 1877 2083 1883
rect 68 1857 83 1863
rect 1085 1857 1123 1863
rect 2029 1857 2067 1863
rect 2221 1857 2252 1863
rect 1544 1837 1596 1843
rect 1544 1806 1550 1814
rect 1558 1806 1564 1814
rect 1572 1806 1578 1814
rect 1586 1806 1592 1814
rect 138 1776 140 1784
rect 698 1776 700 1784
rect 1316 1776 1318 1784
rect 1501 1757 1516 1763
rect 77 1717 115 1723
rect 557 1717 572 1723
rect 589 1717 675 1723
rect 1341 1717 1356 1723
rect 1396 1717 1411 1723
rect 1469 1717 1491 1723
rect 861 1697 876 1703
rect 1460 1636 1462 1644
rect 632 1606 638 1614
rect 646 1606 652 1614
rect 660 1606 666 1614
rect 674 1606 680 1614
rect 557 1577 604 1583
rect 1549 1577 1596 1583
rect 941 1537 956 1543
rect 1412 1517 1427 1523
rect 45 1497 82 1503
rect 2174 1497 2211 1503
rect 509 1477 563 1483
rect 1316 1477 1331 1483
rect 1373 1477 1395 1483
rect 1812 1477 1827 1483
rect 2237 1477 2252 1483
rect 68 1457 83 1463
rect 1544 1406 1550 1414
rect 1558 1406 1564 1414
rect 1572 1406 1578 1414
rect 1586 1406 1592 1414
rect 138 1376 140 1384
rect 852 1376 854 1384
rect 1453 1377 1468 1383
rect 1405 1357 1420 1363
rect 733 1337 748 1343
rect 77 1317 115 1323
rect 637 1317 700 1323
rect 877 1317 915 1323
rect 1837 1277 1852 1283
rect 632 1206 638 1214
rect 646 1206 652 1214
rect 660 1206 666 1214
rect 674 1206 680 1214
rect 1946 1176 1948 1184
rect 148 1137 163 1143
rect 1498 1136 1500 1144
rect 2221 1137 2252 1143
rect 93 1097 108 1103
rect 349 1097 364 1103
rect 1292 1103 1300 1108
rect 1262 1097 1300 1103
rect 1373 1097 1388 1103
rect 1597 1097 1635 1103
rect 157 1077 195 1083
rect 228 1077 243 1083
rect 1597 1083 1603 1097
rect 1725 1097 1763 1103
rect 2077 1103 2083 1123
rect 1949 1097 2003 1103
rect 2013 1097 2067 1103
rect 2077 1097 2092 1103
rect 1517 1077 1603 1083
rect 1764 1077 1779 1083
rect 724 1057 771 1063
rect 2141 1057 2163 1063
rect 1780 1036 1782 1044
rect 1544 1006 1550 1014
rect 1558 1006 1564 1014
rect 1572 1006 1578 1014
rect 1586 1006 1592 1014
rect 621 917 684 923
rect 1117 917 1132 923
rect 1229 897 1244 903
rect 2164 896 2172 904
rect 2188 877 2204 883
rect 516 836 520 844
rect 632 806 638 814
rect 646 806 652 814
rect 660 806 666 814
rect 674 806 680 814
rect 1924 776 1926 784
rect 2234 776 2236 784
rect 2058 736 2060 744
rect 2180 736 2182 744
rect 413 717 428 723
rect 605 717 668 723
rect 1860 716 1868 724
rect 1300 697 1363 703
rect 2205 703 2211 716
rect 2205 697 2227 703
rect 717 677 732 683
rect 1332 677 1347 683
rect 733 657 755 663
rect 1341 657 1356 663
rect 1274 636 1276 644
rect 1544 606 1550 614
rect 1558 606 1564 614
rect 1572 606 1578 614
rect 1586 606 1592 614
rect 456 576 460 584
rect 1924 576 1928 584
rect 381 544 387 563
rect 2180 557 2204 563
rect 205 537 259 543
rect 388 537 403 543
rect 861 537 876 543
rect 637 517 684 523
rect 1101 523 1107 543
rect 1053 517 1091 523
rect 1101 517 1124 523
rect 1116 512 1124 517
rect 1821 523 1827 543
rect 2148 537 2163 543
rect 1821 517 1836 523
rect 1956 517 2019 523
rect 2052 517 2067 523
rect 2173 517 2188 523
rect 2189 497 2195 516
rect 2093 477 2108 483
rect 1044 436 1046 444
rect 632 406 638 414
rect 646 406 652 414
rect 660 406 666 414
rect 674 406 680 414
rect 2106 376 2108 384
rect 829 303 835 323
rect 957 317 972 323
rect 829 297 867 303
rect 877 297 924 303
rect 1204 297 1219 303
rect 1229 297 1266 303
rect 1709 303 1715 323
rect 1709 297 1724 303
rect 1869 303 1875 323
rect 2061 317 2083 323
rect 1789 297 1827 303
rect 1837 297 1875 303
rect 2140 303 2148 308
rect 2125 297 2148 303
rect 1661 277 1676 283
rect 1741 277 1772 283
rect 2125 277 2131 297
rect 2237 297 2252 303
rect 1085 257 1100 263
rect 1636 257 1651 263
rect 1700 256 1708 264
rect 1882 236 1884 244
rect 1544 206 1550 214
rect 1558 206 1564 214
rect 1572 206 1578 214
rect 1586 206 1592 214
rect 1700 157 1715 163
rect 1581 137 1612 143
rect 45 117 82 123
rect 734 117 819 123
rect 900 117 930 123
rect 1404 123 1412 128
rect 1389 117 1412 123
rect 1453 117 1491 123
rect 1501 117 1539 123
rect 1533 97 1539 117
rect 1677 117 1714 123
rect 2132 97 2147 103
rect 2237 77 2252 83
rect 632 6 638 14
rect 646 6 652 14
rect 660 6 666 14
rect 674 6 680 14
<< m2contact >>
rect 638 2006 646 2014
rect 652 2006 660 2014
rect 666 2006 674 2014
rect 364 1976 372 1984
rect 412 1976 420 1984
rect 812 1976 820 1984
rect 860 1976 868 1984
rect 940 1976 948 1984
rect 988 1976 996 1984
rect 1596 1976 1604 1984
rect 1964 1976 1972 1984
rect 2156 1976 2164 1984
rect 1212 1958 1220 1966
rect 1532 1936 1540 1944
rect 364 1916 372 1924
rect 812 1916 820 1924
rect 1212 1912 1220 1920
rect 1500 1916 1508 1924
rect 1964 1916 1972 1924
rect 364 1896 372 1904
rect 812 1896 820 1904
rect 892 1896 900 1904
rect 908 1896 916 1904
rect 956 1896 964 1904
rect 1100 1896 1108 1904
rect 1180 1896 1188 1904
rect 1516 1896 1524 1904
rect 1644 1896 1652 1904
rect 1948 1896 1956 1904
rect 2044 1896 2052 1904
rect 2188 1896 2196 1904
rect 12 1876 20 1884
rect 268 1876 276 1884
rect 716 1876 724 1884
rect 1052 1876 1060 1884
rect 1084 1876 1092 1884
rect 1276 1876 1284 1884
rect 1868 1876 1876 1884
rect 2044 1876 2052 1884
rect 2092 1876 2100 1884
rect 60 1856 68 1864
rect 236 1856 244 1864
rect 684 1856 692 1864
rect 1004 1856 1012 1864
rect 1132 1856 1140 1864
rect 1308 1856 1316 1864
rect 1836 1856 1844 1864
rect 2012 1856 2020 1864
rect 2140 1856 2148 1864
rect 2252 1856 2260 1864
rect 524 1836 532 1844
rect 1468 1836 1476 1844
rect 1596 1836 1604 1844
rect 1676 1836 1684 1844
rect 2204 1836 2212 1844
rect 1550 1806 1558 1814
rect 1564 1806 1572 1814
rect 1578 1806 1586 1814
rect 140 1776 148 1784
rect 700 1776 708 1784
rect 780 1776 788 1784
rect 892 1776 900 1784
rect 1308 1776 1316 1784
rect 2236 1776 2244 1784
rect 60 1756 68 1764
rect 364 1756 372 1764
rect 540 1756 548 1764
rect 572 1756 580 1764
rect 796 1756 804 1764
rect 1052 1756 1060 1764
rect 1388 1756 1396 1764
rect 1420 1756 1428 1764
rect 1436 1756 1444 1764
rect 1516 1756 1524 1764
rect 1580 1756 1588 1764
rect 1740 1756 1748 1764
rect 2076 1756 2084 1764
rect 396 1736 404 1744
rect 764 1736 772 1744
rect 812 1736 820 1744
rect 844 1736 852 1744
rect 1084 1736 1092 1744
rect 1228 1736 1236 1744
rect 1772 1736 1780 1744
rect 2044 1736 2052 1744
rect 44 1716 52 1724
rect 156 1716 164 1724
rect 172 1716 180 1724
rect 396 1716 404 1724
rect 492 1716 500 1724
rect 572 1716 580 1724
rect 716 1716 724 1724
rect 732 1716 740 1724
rect 748 1716 756 1724
rect 828 1716 836 1724
rect 972 1716 980 1724
rect 1180 1716 1188 1724
rect 1260 1716 1268 1724
rect 1276 1716 1284 1724
rect 1292 1716 1300 1724
rect 1356 1716 1364 1724
rect 1388 1716 1396 1724
rect 1660 1716 1668 1724
rect 1884 1716 1892 1724
rect 1948 1716 1956 1724
rect 460 1700 468 1708
rect 876 1696 884 1704
rect 1148 1700 1156 1708
rect 1372 1696 1380 1704
rect 1868 1696 1876 1704
rect 1948 1696 1956 1704
rect 12 1676 20 1684
rect 204 1656 212 1664
rect 1148 1654 1156 1662
rect 460 1636 468 1644
rect 1452 1636 1460 1644
rect 1868 1636 1876 1644
rect 1948 1636 1956 1644
rect 638 1606 646 1614
rect 652 1606 660 1614
rect 666 1606 674 1614
rect 364 1576 372 1584
rect 604 1576 612 1584
rect 652 1576 660 1584
rect 1596 1576 1604 1584
rect 1036 1558 1044 1566
rect 1916 1558 1924 1566
rect 956 1536 964 1544
rect 364 1516 372 1524
rect 412 1516 420 1524
rect 652 1516 660 1524
rect 1036 1512 1044 1520
rect 1324 1516 1332 1524
rect 1404 1516 1412 1524
rect 1916 1512 1924 1520
rect 364 1496 372 1504
rect 444 1496 452 1504
rect 524 1496 532 1504
rect 860 1496 868 1504
rect 1004 1496 1012 1504
rect 1294 1496 1302 1504
rect 1356 1496 1364 1504
rect 1468 1496 1476 1504
rect 1516 1496 1524 1504
rect 1740 1496 1748 1504
rect 1756 1496 1764 1504
rect 1804 1496 1812 1504
rect 1884 1496 1892 1504
rect 1900 1496 1908 1504
rect 12 1476 20 1484
rect 268 1476 276 1484
rect 428 1476 436 1484
rect 460 1476 468 1484
rect 748 1476 756 1484
rect 1100 1476 1108 1484
rect 1308 1476 1316 1484
rect 1452 1476 1460 1484
rect 1612 1476 1620 1484
rect 1772 1476 1780 1484
rect 1804 1476 1812 1484
rect 1980 1476 1988 1484
rect 2252 1476 2260 1484
rect 60 1456 68 1464
rect 236 1456 244 1464
rect 476 1456 484 1464
rect 540 1456 548 1464
rect 780 1456 788 1464
rect 1132 1456 1140 1464
rect 1404 1456 1412 1464
rect 1436 1456 1444 1464
rect 1804 1456 1812 1464
rect 1836 1456 1844 1464
rect 2012 1456 2020 1464
rect 2172 1456 2180 1464
rect 492 1436 500 1444
rect 940 1436 948 1444
rect 1500 1436 1508 1444
rect 1550 1406 1558 1414
rect 1564 1406 1572 1414
rect 1578 1406 1586 1414
rect 140 1376 148 1384
rect 204 1376 212 1384
rect 844 1376 852 1384
rect 956 1376 964 1384
rect 1468 1376 1476 1384
rect 1836 1376 1844 1384
rect 60 1356 68 1364
rect 364 1356 372 1364
rect 588 1356 596 1364
rect 748 1356 756 1364
rect 924 1356 932 1364
rect 1244 1356 1252 1364
rect 1420 1356 1428 1364
rect 1436 1356 1444 1364
rect 1676 1356 1684 1364
rect 2028 1356 2036 1364
rect 396 1336 404 1344
rect 540 1336 548 1344
rect 604 1336 612 1344
rect 748 1336 756 1344
rect 780 1336 788 1344
rect 1068 1336 1076 1344
rect 1212 1336 1220 1344
rect 1644 1336 1652 1344
rect 1996 1336 2004 1344
rect 44 1316 52 1324
rect 156 1316 164 1324
rect 172 1316 180 1324
rect 460 1316 468 1324
rect 556 1316 564 1324
rect 700 1316 708 1324
rect 796 1316 804 1324
rect 812 1316 820 1324
rect 828 1316 836 1324
rect 1116 1316 1124 1324
rect 1756 1316 1764 1324
rect 1900 1316 1908 1324
rect 492 1296 500 1304
rect 588 1296 596 1304
rect 1148 1300 1156 1308
rect 1580 1300 1588 1308
rect 1900 1296 1908 1304
rect 12 1276 20 1284
rect 1852 1276 1860 1284
rect 1756 1254 1764 1262
rect 492 1236 500 1244
rect 748 1236 756 1244
rect 1148 1236 1156 1244
rect 1900 1236 1908 1244
rect 2188 1236 2196 1244
rect 638 1206 646 1214
rect 652 1206 660 1214
rect 666 1206 674 1214
rect 124 1176 132 1184
rect 668 1176 676 1184
rect 780 1176 788 1184
rect 972 1176 980 1184
rect 1260 1176 1268 1184
rect 1340 1176 1348 1184
rect 1436 1176 1444 1184
rect 1948 1176 1956 1184
rect 1836 1156 1844 1164
rect 12 1136 20 1144
rect 140 1136 148 1144
rect 1324 1136 1332 1144
rect 1500 1136 1508 1144
rect 1900 1136 1908 1144
rect 2252 1136 2260 1144
rect 284 1116 292 1124
rect 668 1116 676 1124
rect 972 1116 980 1124
rect 1404 1116 1412 1124
rect 1468 1116 1476 1124
rect 1740 1116 1748 1124
rect 1916 1116 1924 1124
rect 1980 1116 1988 1124
rect 44 1096 52 1104
rect 108 1096 116 1104
rect 172 1096 180 1104
rect 252 1096 260 1104
rect 300 1096 308 1104
rect 364 1096 372 1104
rect 460 1096 468 1104
rect 668 1096 676 1104
rect 988 1096 996 1104
rect 1004 1096 1012 1104
rect 1308 1096 1316 1104
rect 1388 1096 1396 1104
rect 1420 1096 1428 1104
rect 1500 1096 1508 1104
rect 1564 1096 1572 1104
rect 60 1076 68 1084
rect 220 1076 228 1084
rect 268 1076 276 1084
rect 316 1076 324 1084
rect 378 1076 386 1084
rect 572 1076 580 1084
rect 796 1076 804 1084
rect 924 1076 932 1084
rect 1068 1076 1076 1084
rect 1708 1096 1716 1104
rect 1820 1096 1828 1104
rect 1868 1096 1876 1104
rect 2092 1096 2100 1104
rect 2188 1096 2196 1104
rect 1644 1076 1652 1084
rect 1692 1076 1700 1084
rect 1756 1076 1764 1084
rect 1804 1076 1812 1084
rect 1964 1076 1972 1084
rect 2028 1076 2036 1084
rect 2044 1076 2052 1084
rect 2108 1076 2116 1084
rect 108 1056 116 1064
rect 140 1056 148 1064
rect 220 1056 228 1064
rect 348 1056 356 1064
rect 540 1056 548 1064
rect 716 1056 724 1064
rect 1100 1056 1108 1064
rect 1356 1056 1364 1064
rect 1388 1056 1396 1064
rect 1452 1056 1460 1064
rect 1532 1056 1540 1064
rect 1676 1056 1684 1064
rect 1852 1056 1860 1064
rect 2172 1056 2180 1064
rect 204 1036 212 1044
rect 1660 1036 1668 1044
rect 1772 1036 1780 1044
rect 2076 1036 2084 1044
rect 2124 1036 2132 1044
rect 1550 1006 1558 1014
rect 1564 1006 1572 1014
rect 1578 1006 1586 1014
rect 28 976 36 984
rect 412 976 420 984
rect 1084 976 1092 984
rect 1356 976 1364 984
rect 2092 976 2100 984
rect 188 956 196 964
rect 700 956 708 964
rect 860 956 868 964
rect 1324 956 1332 964
rect 1516 956 1524 964
rect 1900 956 1908 964
rect 220 936 228 944
rect 364 936 372 944
rect 460 936 468 944
rect 476 936 484 944
rect 572 936 580 944
rect 588 936 596 944
rect 892 936 900 944
rect 1548 936 1556 944
rect 1868 936 1876 944
rect 2124 936 2132 944
rect 2140 936 2148 944
rect 300 916 308 924
rect 396 916 404 924
rect 444 916 452 924
rect 684 916 692 924
rect 988 916 996 924
rect 1068 916 1076 924
rect 1132 916 1140 924
rect 1212 916 1220 924
rect 1260 916 1268 924
rect 1308 916 1316 924
rect 1436 916 1444 924
rect 1612 916 1620 924
rect 1772 916 1780 924
rect 2156 916 2164 924
rect 2220 916 2228 924
rect 316 896 324 904
rect 412 896 420 904
rect 988 896 996 904
rect 1244 896 1252 904
rect 1644 896 1652 904
rect 1804 900 1812 908
rect 2092 896 2100 904
rect 2156 896 2164 904
rect 2204 896 2212 904
rect 1164 876 1172 884
rect 1196 876 1204 884
rect 1276 876 1284 884
rect 2204 876 2212 884
rect 2236 876 2244 884
rect 1804 854 1812 862
rect 2220 856 2228 864
rect 28 836 36 844
rect 316 836 324 844
rect 508 836 516 844
rect 988 836 996 844
rect 1036 836 1044 844
rect 1180 836 1188 844
rect 1260 836 1268 844
rect 1356 836 1364 844
rect 1644 836 1652 844
rect 2060 836 2068 844
rect 638 806 646 814
rect 652 806 660 814
rect 666 806 674 814
rect 316 776 324 784
rect 684 776 692 784
rect 1180 776 1188 784
rect 1196 776 1204 784
rect 1516 776 1524 784
rect 1916 776 1924 784
rect 2236 776 2244 784
rect 876 758 884 766
rect 2108 756 2116 764
rect 412 736 420 744
rect 2060 736 2068 744
rect 2124 736 2132 744
rect 2172 736 2180 744
rect 316 716 324 724
rect 428 716 436 724
rect 540 716 548 724
rect 668 716 676 724
rect 748 716 756 724
rect 876 712 884 720
rect 1516 716 1524 724
rect 1852 716 1860 724
rect 1884 716 1892 724
rect 1948 716 1956 724
rect 2028 716 2036 724
rect 2092 716 2100 724
rect 2204 716 2212 724
rect 300 696 308 704
rect 316 696 324 704
rect 380 696 388 704
rect 460 696 468 704
rect 492 696 500 704
rect 572 696 580 704
rect 700 696 708 704
rect 780 696 788 704
rect 828 696 836 704
rect 1052 696 1060 704
rect 1134 696 1142 704
rect 1228 696 1236 704
rect 1292 696 1300 704
rect 1516 696 1524 704
rect 1612 696 1620 704
rect 1852 696 1860 704
rect 1916 696 1924 704
rect 1980 696 1988 704
rect 2012 696 2020 704
rect 2060 696 2068 704
rect 2108 696 2116 704
rect 2172 696 2180 704
rect 220 676 228 684
rect 364 676 372 684
rect 476 676 484 684
rect 508 676 516 684
rect 556 676 564 684
rect 588 676 596 684
rect 732 676 740 684
rect 796 676 804 684
rect 940 676 948 684
rect 1244 676 1252 684
rect 1276 676 1284 684
rect 1324 676 1332 684
rect 1612 676 1620 684
rect 1836 676 1844 684
rect 1900 676 1908 684
rect 1996 676 2004 684
rect 2076 676 2084 684
rect 2156 676 2164 684
rect 188 656 196 664
rect 540 656 548 664
rect 668 656 676 664
rect 972 656 980 664
rect 1164 656 1172 664
rect 1212 656 1220 664
rect 1356 656 1364 664
rect 1644 656 1652 664
rect 1964 656 1972 664
rect 2252 656 2260 664
rect 28 636 36 644
rect 412 636 420 644
rect 428 636 436 644
rect 684 636 692 644
rect 1276 636 1284 644
rect 1340 636 1348 644
rect 1804 636 1812 644
rect 1550 606 1558 614
rect 1564 606 1572 614
rect 1578 606 1586 614
rect 268 576 276 584
rect 460 576 468 584
rect 748 576 756 584
rect 1036 576 1044 584
rect 1260 576 1268 584
rect 1756 576 1764 584
rect 1916 576 1924 584
rect 2124 576 2132 584
rect 2188 576 2196 584
rect 220 556 228 564
rect 284 556 292 564
rect 348 556 356 564
rect 364 556 372 564
rect 716 556 724 564
rect 1020 556 1028 564
rect 1420 556 1428 564
rect 1868 556 1876 564
rect 2108 556 2116 564
rect 2140 556 2148 564
rect 2172 556 2180 564
rect 12 536 20 544
rect 316 536 324 544
rect 380 536 388 544
rect 492 536 500 544
rect 876 536 884 544
rect 1004 536 1012 544
rect 44 516 52 524
rect 92 516 100 524
rect 124 516 132 524
rect 172 516 180 524
rect 188 516 196 524
rect 236 516 244 524
rect 300 516 308 524
rect 508 516 516 524
rect 524 516 532 524
rect 572 516 580 524
rect 684 516 692 524
rect 700 516 708 524
rect 1452 536 1460 544
rect 1644 536 1652 544
rect 1676 536 1684 544
rect 1708 536 1716 544
rect 1772 536 1780 544
rect 1132 516 1140 524
rect 1212 516 1220 524
rect 1516 516 1524 524
rect 1660 516 1668 524
rect 1724 516 1732 524
rect 1804 516 1812 524
rect 1884 536 1892 544
rect 1980 536 1988 544
rect 2044 536 2052 544
rect 2140 536 2148 544
rect 2220 536 2228 544
rect 1836 516 1844 524
rect 1948 516 1956 524
rect 2028 516 2036 524
rect 2044 516 2052 524
rect 2188 516 2196 524
rect 204 496 212 504
rect 1068 496 1076 504
rect 1116 496 1124 504
rect 1228 496 1236 504
rect 1548 496 1556 504
rect 1692 496 1700 504
rect 1772 496 1780 504
rect 1996 496 2004 504
rect 60 476 68 484
rect 604 476 612 484
rect 1148 476 1156 484
rect 1196 476 1204 484
rect 1836 476 1844 484
rect 2108 476 2116 484
rect 1212 456 1220 464
rect 140 436 148 444
rect 348 436 356 444
rect 556 436 564 444
rect 748 436 756 444
rect 1036 436 1044 444
rect 1132 436 1140 444
rect 1548 436 1556 444
rect 638 406 646 414
rect 652 406 660 414
rect 666 406 674 414
rect 28 376 36 384
rect 60 376 68 384
rect 348 376 356 384
rect 1548 376 1556 384
rect 2108 376 2116 384
rect 2236 376 2244 384
rect 460 358 468 366
rect 1052 356 1060 364
rect 1932 356 1940 364
rect 2156 356 2164 364
rect 716 336 724 344
rect 844 336 852 344
rect 1036 336 1044 344
rect 1084 336 1092 344
rect 1948 336 1956 344
rect 2172 336 2180 344
rect 348 316 356 324
rect 460 312 468 320
rect 332 296 340 304
rect 348 296 356 304
rect 444 296 452 304
rect 636 296 644 304
rect 972 316 980 324
rect 1004 316 1012 324
rect 1116 316 1124 324
rect 1548 316 1556 324
rect 924 296 932 304
rect 988 296 996 304
rect 1020 296 1028 304
rect 1100 296 1108 304
rect 1164 296 1172 304
rect 1196 296 1204 304
rect 1340 296 1348 304
rect 1516 296 1524 304
rect 1852 316 1860 324
rect 1724 296 1732 304
rect 1916 316 1924 324
rect 1980 316 1988 324
rect 2140 316 2148 324
rect 1932 296 1940 304
rect 2012 296 2020 304
rect 2108 296 2116 304
rect 252 276 260 284
rect 524 276 532 284
rect 796 276 804 284
rect 812 276 820 284
rect 892 276 900 284
rect 908 276 916 284
rect 956 276 964 284
rect 1180 276 1188 284
rect 1452 276 1460 284
rect 1676 276 1684 284
rect 1772 276 1780 284
rect 1804 276 1812 284
rect 1900 276 1908 284
rect 1996 276 2004 284
rect 2028 276 2036 284
rect 2156 296 2164 304
rect 2252 296 2260 304
rect 12 256 20 264
rect 220 256 228 264
rect 556 256 564 264
rect 972 256 980 264
rect 1100 256 1108 264
rect 1196 256 1204 264
rect 1420 256 1428 264
rect 1628 256 1636 264
rect 1708 256 1716 264
rect 1756 256 1764 264
rect 1772 256 1780 264
rect 2044 256 2052 264
rect 2204 256 2212 264
rect 1132 236 1140 244
rect 1260 236 1268 244
rect 1884 236 1892 244
rect 1550 206 1558 214
rect 1564 206 1572 214
rect 1578 206 1586 214
rect 76 176 84 184
rect 732 176 740 184
rect 1372 176 1380 184
rect 2092 176 2100 184
rect 2108 176 2116 184
rect 2172 176 2180 184
rect 236 156 244 164
rect 572 156 580 164
rect 1084 156 1092 164
rect 1356 156 1364 164
rect 1532 156 1540 164
rect 1692 156 1700 164
rect 1868 156 1876 164
rect 2124 156 2132 164
rect 2156 156 2164 164
rect 2188 156 2196 164
rect 268 136 276 144
rect 540 136 548 144
rect 1116 136 1124 144
rect 1404 136 1412 144
rect 1468 136 1476 144
rect 1612 136 1620 144
rect 1900 136 1908 144
rect 2044 136 2052 144
rect 348 116 356 124
rect 364 116 372 124
rect 444 116 452 124
rect 892 116 900 124
rect 1212 116 1220 124
rect 1260 116 1268 124
rect 1308 116 1316 124
rect 1420 116 1428 124
rect 364 96 372 104
rect 444 96 452 104
rect 1212 96 1220 104
rect 1516 96 1524 104
rect 1564 116 1572 124
rect 1788 116 1796 124
rect 2060 116 2068 124
rect 2204 116 2212 124
rect 1996 96 2004 104
rect 2092 96 2100 104
rect 2124 96 2132 104
rect 12 76 20 84
rect 2252 76 2260 84
rect 364 36 372 44
rect 444 36 452 44
rect 844 36 852 44
rect 860 36 868 44
rect 1212 36 1220 44
rect 1292 36 1300 44
rect 1340 36 1348 44
rect 1644 36 1652 44
rect 1996 36 2004 44
rect 638 6 646 14
rect 652 6 660 14
rect 666 6 674 14
<< metal2 >>
rect 413 2037 435 2043
rect 413 1984 419 2037
rect 632 2006 638 2014
rect 646 2006 652 2014
rect 660 2006 666 2014
rect 674 2006 680 2014
rect 861 1984 867 2043
rect 925 2037 947 2043
rect 973 2037 995 2043
rect 1373 2037 1395 2043
rect 941 1984 947 2037
rect 989 1984 995 2037
rect 365 1924 371 1976
rect 813 1924 819 1976
rect 1213 1920 1219 1958
rect 13 1884 19 1896
rect 61 1764 67 1856
rect 141 1784 147 1876
rect 173 1724 179 1816
rect 237 1764 243 1856
rect 365 1804 371 1896
rect 13 1684 19 1696
rect 45 1664 51 1716
rect 13 1484 19 1496
rect 45 1324 51 1376
rect 61 1364 67 1456
rect 141 1384 147 1476
rect 157 1343 163 1716
rect 173 1604 179 1716
rect 237 1464 243 1756
rect 397 1744 403 1776
rect 493 1724 499 1796
rect 573 1764 579 1836
rect 685 1764 691 1856
rect 717 1823 723 1876
rect 701 1817 723 1823
rect 701 1784 707 1817
rect 365 1524 371 1576
rect 397 1504 403 1716
rect 461 1644 467 1700
rect 541 1664 547 1756
rect 733 1724 739 1816
rect 813 1804 819 1896
rect 893 1784 899 1896
rect 909 1884 915 1896
rect 845 1744 851 1756
rect 909 1744 915 1876
rect 413 1484 419 1516
rect 429 1464 435 1476
rect 365 1364 371 1456
rect 141 1337 163 1343
rect 13 1284 19 1296
rect 125 1184 131 1216
rect 141 1144 147 1337
rect 157 1224 163 1316
rect 285 1124 291 1276
rect 365 1244 371 1356
rect 493 1344 499 1436
rect 525 1324 531 1496
rect 541 1484 547 1656
rect 605 1584 611 1676
rect 632 1606 638 1614
rect 646 1606 652 1614
rect 660 1606 666 1614
rect 674 1606 680 1614
rect 653 1524 659 1576
rect 749 1504 755 1716
rect 541 1384 547 1456
rect 749 1424 755 1476
rect 781 1423 787 1456
rect 765 1417 787 1423
rect 541 1344 547 1376
rect 605 1324 611 1336
rect 173 1104 179 1116
rect 253 1104 259 1116
rect 45 1064 51 1096
rect 61 1084 67 1096
rect 109 1084 115 1096
rect 109 1064 115 1076
rect 269 1064 275 1076
rect 29 1057 44 1063
rect 29 984 35 1057
rect 205 1003 211 1036
rect 205 997 227 1003
rect 29 684 35 836
rect 189 664 195 956
rect 221 944 227 997
rect 285 944 291 1116
rect 301 1064 307 1096
rect 317 1084 323 1216
rect 461 1104 467 1316
rect 493 1244 499 1296
rect 589 1284 595 1296
rect 349 1044 355 1056
rect 381 984 387 1076
rect 541 1064 547 1236
rect 632 1206 638 1214
rect 646 1206 652 1214
rect 660 1206 666 1214
rect 674 1206 680 1214
rect 669 1124 675 1176
rect 573 1084 579 1096
rect 413 984 419 1036
rect 301 704 307 916
rect 365 904 371 936
rect 397 924 403 956
rect 413 904 419 936
rect 445 924 451 1056
rect 701 983 707 1316
rect 685 977 707 983
rect 477 944 483 976
rect 589 924 595 936
rect 685 924 691 977
rect 717 963 723 1056
rect 708 957 723 963
rect 701 944 707 956
rect 749 944 755 1236
rect 765 1064 771 1417
rect 845 1384 851 1416
rect 781 1324 787 1336
rect 797 1324 803 1336
rect 813 1324 819 1336
rect 781 1184 787 1316
rect 797 1144 803 1316
rect 877 1284 883 1696
rect 797 1064 803 1076
rect 909 1024 915 1736
rect 957 1544 963 1896
rect 1005 1864 1011 1896
rect 1053 1824 1059 1876
rect 973 1724 979 1796
rect 1053 1764 1059 1796
rect 973 1504 979 1716
rect 1053 1624 1059 1756
rect 1085 1744 1091 1876
rect 1101 1824 1107 1896
rect 1133 1864 1139 1876
rect 1181 1724 1187 1896
rect 1277 1784 1283 1876
rect 1309 1804 1315 1856
rect 1229 1724 1235 1736
rect 1341 1724 1347 1816
rect 1389 1764 1395 2037
rect 1597 1984 1603 2043
rect 1421 1764 1427 1776
rect 1261 1704 1267 1716
rect 1149 1662 1155 1700
rect 1293 1684 1299 1716
rect 1037 1520 1043 1558
rect 925 1437 940 1443
rect 925 1364 931 1437
rect 957 1384 963 1456
rect 1005 1324 1011 1496
rect 1133 1464 1139 1616
rect 925 1084 931 1296
rect 973 1124 979 1176
rect 1005 1104 1011 1316
rect 1069 1304 1075 1336
rect 317 844 323 896
rect 317 724 323 776
rect 413 744 419 896
rect 429 724 435 736
rect 461 704 467 916
rect 685 843 691 916
rect 685 837 707 843
rect 324 697 339 703
rect 29 563 35 636
rect 189 584 195 656
rect 221 624 227 676
rect 221 564 227 596
rect 269 584 275 616
rect 285 564 291 616
rect 29 557 44 563
rect 45 524 51 556
rect 317 544 323 556
rect 93 524 99 536
rect 29 384 35 516
rect 61 484 67 496
rect 93 384 99 516
rect 173 504 179 516
rect 237 484 243 516
rect 301 484 307 516
rect 13 184 19 256
rect 141 144 147 436
rect 221 264 227 316
rect 253 284 259 396
rect 333 304 339 697
rect 509 684 515 836
rect 632 806 638 814
rect 646 806 652 814
rect 660 806 666 814
rect 674 806 680 814
rect 701 783 707 837
rect 692 777 707 783
rect 749 724 755 736
rect 756 717 771 723
rect 557 684 563 696
rect 573 684 579 696
rect 484 677 499 683
rect 365 604 371 676
rect 413 584 419 636
rect 429 624 435 636
rect 461 584 467 636
rect 349 564 355 576
rect 493 544 499 677
rect 557 644 563 676
rect 589 664 595 676
rect 669 664 675 716
rect 701 704 707 716
rect 525 524 531 556
rect 685 524 691 636
rect 749 584 755 636
rect 349 404 355 436
rect 349 324 355 376
rect 461 320 467 358
rect 557 344 563 436
rect 632 406 638 414
rect 646 406 652 414
rect 660 406 666 414
rect 674 406 680 414
rect 717 363 723 556
rect 717 357 739 363
rect 221 203 227 256
rect 221 197 243 203
rect 237 164 243 197
rect 349 124 355 296
rect 445 124 451 296
rect 557 264 563 316
rect 557 203 563 256
rect 557 197 579 203
rect 573 164 579 197
rect 733 184 739 357
rect 749 324 755 436
rect 765 324 771 717
rect 781 704 787 1016
rect 925 1004 931 1076
rect 989 984 995 1096
rect 989 924 995 976
rect 1069 963 1075 1076
rect 1101 1064 1107 1456
rect 1245 1364 1251 1456
rect 1149 1244 1155 1300
rect 1213 1244 1219 1336
rect 1261 1184 1267 1236
rect 1341 1184 1347 1716
rect 1453 1703 1459 1916
rect 1469 1784 1475 1836
rect 1437 1697 1459 1703
rect 1357 1484 1363 1496
rect 1405 1464 1411 1496
rect 1437 1464 1443 1697
rect 1453 1484 1459 1636
rect 1437 1383 1443 1456
rect 1469 1384 1475 1476
rect 1421 1377 1443 1383
rect 1421 1364 1427 1377
rect 1437 1244 1443 1356
rect 1101 964 1107 1056
rect 1069 957 1091 963
rect 1069 924 1075 936
rect 989 844 995 896
rect 1037 803 1043 836
rect 1085 804 1091 957
rect 1133 924 1139 936
rect 1245 904 1251 1176
rect 1309 1104 1315 1156
rect 1469 1124 1475 1156
rect 1485 1144 1491 1896
rect 1533 1864 1539 1936
rect 1501 1484 1507 1856
rect 1604 1837 1619 1843
rect 1517 1764 1523 1836
rect 1544 1806 1550 1814
rect 1558 1806 1564 1814
rect 1572 1806 1578 1814
rect 1586 1806 1592 1814
rect 1517 1504 1523 1696
rect 1597 1584 1603 1716
rect 1613 1504 1619 1837
rect 1629 1483 1635 2043
rect 1821 2004 1827 2043
rect 2013 2037 2035 2043
rect 2157 2037 2179 2043
rect 1645 1784 1651 1896
rect 1869 1884 1875 1996
rect 1965 1924 1971 1976
rect 1677 1804 1683 1836
rect 1741 1504 1747 1756
rect 1773 1744 1779 1796
rect 1837 1764 1843 1856
rect 1949 1724 1955 1896
rect 2013 1864 2019 2037
rect 2157 1984 2163 2037
rect 2045 1744 2051 1876
rect 2141 1864 2147 1896
rect 1869 1644 1875 1696
rect 1885 1504 1891 1716
rect 1949 1644 1955 1696
rect 1917 1520 1923 1558
rect 1620 1477 1635 1483
rect 1501 1344 1507 1436
rect 1544 1406 1550 1414
rect 1558 1406 1564 1414
rect 1572 1406 1578 1414
rect 1586 1406 1592 1414
rect 1741 1404 1747 1496
rect 1805 1444 1811 1456
rect 1677 1364 1683 1396
rect 1837 1384 1843 1436
rect 1901 1324 1907 1496
rect 1981 1484 1987 1496
rect 2013 1404 2019 1456
rect 2020 1397 2035 1403
rect 2029 1364 2035 1397
rect 1581 1308 1587 1316
rect 1757 1262 1763 1316
rect 1165 884 1171 896
rect 1277 884 1283 1096
rect 1453 1064 1459 1116
rect 1325 964 1331 1056
rect 1357 1044 1363 1056
rect 1357 984 1363 996
rect 1181 824 1187 836
rect 1037 797 1059 803
rect 877 720 883 758
rect 1053 704 1059 797
rect 1181 784 1187 796
rect 1197 784 1203 876
rect 1261 703 1267 836
rect 1261 697 1283 703
rect 797 664 803 676
rect 797 344 803 656
rect 797 284 803 316
rect 829 304 835 696
rect 1213 664 1219 676
rect 973 644 979 656
rect 877 544 883 596
rect 1037 584 1043 616
rect 909 284 915 476
rect 1005 364 1011 416
rect 925 304 931 336
rect 1005 324 1011 356
rect 1037 344 1043 436
rect 1085 344 1091 356
rect 1101 323 1107 536
rect 1117 504 1123 516
rect 1133 504 1139 516
rect 1133 344 1139 436
rect 1165 364 1171 656
rect 1213 504 1219 516
rect 1229 504 1235 696
rect 1277 684 1283 697
rect 1293 684 1299 696
rect 1325 684 1331 956
rect 1389 924 1395 1056
rect 1453 1004 1459 1056
rect 1565 1044 1571 1096
rect 1645 1084 1651 1176
rect 1853 1104 1859 1276
rect 1901 1244 1907 1296
rect 1997 1224 2003 1336
rect 1949 1184 1955 1216
rect 1901 1124 1907 1136
rect 1917 1124 1923 1136
rect 1869 1104 1875 1116
rect 1981 1104 1987 1116
rect 1709 1063 1715 1096
rect 1709 1057 1731 1063
rect 1544 1006 1550 1014
rect 1558 1006 1564 1014
rect 1572 1006 1578 1014
rect 1586 1006 1592 1014
rect 1437 904 1443 916
rect 1517 843 1523 956
rect 1517 837 1539 843
rect 1245 624 1251 676
rect 1261 584 1267 676
rect 1277 524 1283 636
rect 1197 484 1203 496
rect 1085 317 1107 323
rect 893 264 899 276
rect 893 124 899 256
rect 909 144 915 276
rect 973 264 979 316
rect 1085 164 1091 317
rect 1101 284 1107 296
rect 1117 284 1123 316
rect 1165 304 1171 336
rect 1197 304 1203 476
rect 1229 424 1235 496
rect 1181 264 1187 276
rect 1133 203 1139 236
rect 1117 197 1139 203
rect 1117 144 1123 197
rect 1261 184 1267 236
rect 1293 164 1299 676
rect 1357 664 1363 836
rect 1517 724 1523 776
rect 1341 484 1347 636
rect 1421 564 1427 636
rect 1421 544 1427 556
rect 1261 124 1267 156
rect 1309 124 1315 176
rect 1341 124 1347 296
rect 1421 264 1427 536
rect 1517 524 1523 696
rect 1533 644 1539 837
rect 1613 704 1619 916
rect 1645 844 1651 896
rect 1645 644 1651 656
rect 1544 606 1550 614
rect 1558 606 1564 614
rect 1572 606 1578 614
rect 1586 606 1592 614
rect 1645 544 1651 576
rect 1725 524 1731 1057
rect 1757 1044 1763 1076
rect 1773 944 1779 1036
rect 1805 1024 1811 1076
rect 1853 1064 1859 1096
rect 1965 1044 1971 1076
rect 1805 862 1811 900
rect 1869 844 1875 936
rect 1917 784 1923 836
rect 1885 724 1891 756
rect 1949 724 1955 736
rect 1981 724 1987 1096
rect 2029 964 2035 1076
rect 2045 1064 2051 1076
rect 2109 1064 2115 1076
rect 2077 924 2083 1036
rect 2093 984 2099 1016
rect 2141 944 2147 956
rect 2157 944 2163 1856
rect 2189 1104 2195 1236
rect 2189 1084 2195 1096
rect 2173 964 2179 1056
rect 2061 804 2067 836
rect 1757 584 1763 696
rect 1901 684 1907 716
rect 2029 704 2035 716
rect 2077 704 2083 916
rect 2125 884 2131 936
rect 2173 824 2179 916
rect 2189 903 2195 1056
rect 2205 944 2211 1836
rect 2237 1784 2243 1896
rect 2253 1484 2259 1496
rect 2221 924 2227 1096
rect 2189 897 2204 903
rect 1837 524 1843 536
rect 1517 304 1523 516
rect 1549 444 1555 496
rect 1693 444 1699 496
rect 1725 464 1731 516
rect 1773 504 1779 516
rect 1805 484 1811 516
rect 1549 324 1555 376
rect 1421 244 1427 256
rect 1357 164 1363 176
rect 1453 164 1459 276
rect 1357 124 1363 156
rect 1469 144 1475 176
rect 1517 124 1523 296
rect 1544 206 1550 214
rect 1558 206 1564 214
rect 1572 206 1578 214
rect 1586 206 1592 214
rect 1613 204 1619 276
rect 1565 124 1571 176
rect 1613 144 1619 196
rect 1693 164 1699 256
rect 1725 144 1731 296
rect 1757 264 1763 276
rect 1821 224 1827 516
rect 1837 484 1843 496
rect 1853 324 1859 656
rect 1869 564 1875 636
rect 1901 584 1907 676
rect 1917 584 1923 696
rect 2013 664 2019 696
rect 2061 664 2067 696
rect 2125 664 2131 696
rect 1869 524 1875 556
rect 1885 484 1891 536
rect 1853 204 1859 316
rect 1885 264 1891 476
rect 1949 364 1955 516
rect 1997 504 2003 576
rect 2029 524 2035 656
rect 2125 584 2131 656
rect 2141 564 2147 576
rect 2125 557 2140 563
rect 1901 284 1907 356
rect 1933 344 1939 356
rect 1997 323 2003 496
rect 2109 484 2115 496
rect 2109 384 2115 436
rect 1988 317 2003 323
rect 1933 244 1939 296
rect 1997 264 2003 276
rect 1869 164 1875 236
rect 1885 203 1891 236
rect 1885 197 1907 203
rect 1901 144 1907 197
rect 2029 143 2035 276
rect 2061 164 2067 296
rect 2093 184 2099 236
rect 2125 164 2131 557
rect 2157 383 2163 636
rect 2189 584 2195 897
rect 2205 864 2211 876
rect 2221 864 2227 876
rect 2237 843 2243 876
rect 2221 837 2243 843
rect 2221 763 2227 837
rect 2237 784 2243 816
rect 2221 757 2243 763
rect 2221 544 2227 576
rect 2189 524 2195 536
rect 2237 384 2243 757
rect 2253 664 2259 676
rect 2141 377 2163 383
rect 2141 324 2147 377
rect 2157 344 2163 356
rect 2173 304 2179 336
rect 2253 304 2259 336
rect 2157 264 2163 296
rect 2157 164 2163 256
rect 2173 184 2179 296
rect 2029 137 2044 143
rect 1613 104 1619 136
rect 2061 124 2067 156
rect 2205 124 2211 216
rect 13 84 19 96
rect 365 44 371 96
rect 445 44 451 96
rect 1213 44 1219 96
rect 1997 44 2003 96
rect 2253 84 2259 96
rect 845 24 851 36
rect 632 6 638 14
rect 646 6 652 14
rect 660 6 666 14
rect 674 6 680 14
rect 813 -23 819 16
rect 861 -17 867 36
rect 1293 -17 1299 36
rect 1341 -17 1347 36
rect 861 -23 883 -17
rect 1277 -23 1299 -17
rect 1325 -23 1347 -17
rect 1645 -17 1651 36
rect 1645 -23 1667 -17
<< m3contact >>
rect 638 2006 646 2014
rect 652 2006 660 2014
rect 666 2006 674 2014
rect 12 1896 20 1904
rect 892 1896 900 1904
rect 1004 1896 1012 1904
rect 140 1876 148 1884
rect 268 1876 276 1884
rect 172 1816 180 1824
rect 524 1836 532 1844
rect 572 1836 580 1844
rect 364 1796 372 1804
rect 492 1796 500 1804
rect 396 1776 404 1784
rect 236 1756 244 1764
rect 364 1756 372 1764
rect 12 1696 20 1704
rect 44 1656 52 1664
rect 12 1496 20 1504
rect 140 1476 148 1484
rect 44 1376 52 1384
rect 204 1656 212 1664
rect 172 1596 180 1604
rect 732 1816 740 1824
rect 684 1756 692 1764
rect 812 1796 820 1804
rect 908 1876 916 1884
rect 780 1776 788 1784
rect 796 1756 804 1764
rect 844 1756 852 1764
rect 764 1736 772 1744
rect 812 1736 820 1744
rect 908 1736 916 1744
rect 572 1716 580 1724
rect 716 1716 724 1724
rect 748 1716 756 1724
rect 828 1716 836 1724
rect 604 1676 612 1684
rect 540 1656 548 1664
rect 364 1496 372 1504
rect 396 1496 404 1504
rect 444 1496 452 1504
rect 524 1496 532 1504
rect 268 1476 276 1484
rect 412 1476 420 1484
rect 460 1476 468 1484
rect 236 1456 244 1464
rect 364 1456 372 1464
rect 428 1456 436 1464
rect 476 1456 484 1464
rect 204 1376 212 1384
rect 12 1296 20 1304
rect 124 1216 132 1224
rect 172 1316 180 1324
rect 284 1276 292 1284
rect 156 1216 164 1224
rect 12 1136 20 1144
rect 396 1336 404 1344
rect 492 1336 500 1344
rect 638 1606 646 1614
rect 652 1606 660 1614
rect 666 1606 674 1614
rect 748 1496 756 1504
rect 860 1496 868 1504
rect 540 1476 548 1484
rect 748 1416 756 1424
rect 540 1376 548 1384
rect 588 1356 596 1364
rect 748 1356 756 1364
rect 748 1336 756 1344
rect 524 1316 532 1324
rect 556 1316 564 1324
rect 604 1316 612 1324
rect 364 1236 372 1244
rect 316 1216 324 1224
rect 172 1116 180 1124
rect 252 1116 260 1124
rect 60 1096 68 1104
rect 108 1076 116 1084
rect 220 1076 228 1084
rect 44 1056 52 1064
rect 140 1056 148 1064
rect 220 1056 228 1064
rect 268 1056 276 1064
rect 28 676 36 684
rect 588 1276 596 1284
rect 540 1236 548 1244
rect 364 1096 372 1104
rect 380 1076 386 1084
rect 386 1076 388 1084
rect 300 1056 308 1064
rect 348 1036 356 1044
rect 638 1206 646 1214
rect 652 1206 660 1214
rect 666 1206 674 1214
rect 572 1096 580 1104
rect 668 1096 676 1104
rect 444 1056 452 1064
rect 540 1056 548 1064
rect 412 1036 420 1044
rect 380 976 388 984
rect 396 956 404 964
rect 284 936 292 944
rect 412 936 420 944
rect 476 976 484 984
rect 460 936 468 944
rect 572 936 580 944
rect 844 1416 852 1424
rect 796 1336 804 1344
rect 812 1336 820 1344
rect 780 1316 788 1324
rect 828 1316 836 1324
rect 876 1276 884 1284
rect 796 1136 804 1144
rect 764 1056 772 1064
rect 796 1056 804 1064
rect 1052 1816 1060 1824
rect 972 1796 980 1804
rect 1052 1796 1060 1804
rect 1132 1876 1140 1884
rect 1100 1816 1108 1824
rect 1340 1816 1348 1824
rect 1308 1796 1316 1804
rect 1276 1776 1284 1784
rect 1308 1776 1316 1784
rect 1452 1916 1460 1924
rect 1500 1916 1508 1924
rect 1420 1776 1428 1784
rect 1436 1756 1444 1764
rect 1180 1716 1188 1724
rect 1228 1716 1236 1724
rect 1276 1716 1284 1724
rect 1340 1716 1348 1724
rect 1356 1716 1364 1724
rect 1388 1716 1396 1724
rect 1260 1696 1268 1704
rect 1292 1676 1300 1684
rect 1052 1616 1060 1624
rect 1132 1616 1140 1624
rect 972 1496 980 1504
rect 956 1456 964 1464
rect 1100 1476 1108 1484
rect 1324 1516 1332 1524
rect 1292 1496 1294 1504
rect 1294 1496 1300 1504
rect 1308 1476 1316 1484
rect 1100 1456 1108 1464
rect 1132 1456 1140 1464
rect 1244 1456 1252 1464
rect 1004 1316 1012 1324
rect 924 1296 932 1304
rect 1068 1296 1076 1304
rect 988 1096 996 1104
rect 780 1016 788 1024
rect 908 1016 916 1024
rect 700 936 708 944
rect 748 936 756 944
rect 444 916 452 924
rect 460 916 468 924
rect 588 916 596 924
rect 364 896 372 904
rect 428 736 436 744
rect 220 616 228 624
rect 268 616 276 624
rect 284 616 292 624
rect 220 596 228 604
rect 188 576 196 584
rect 44 556 52 564
rect 220 556 228 564
rect 316 556 324 564
rect 12 536 20 544
rect 92 536 100 544
rect 28 516 36 524
rect 124 516 132 524
rect 188 516 196 524
rect 60 496 68 504
rect 172 496 180 504
rect 204 496 212 504
rect 236 476 244 484
rect 300 476 308 484
rect 60 376 68 384
rect 92 376 100 384
rect 12 176 20 184
rect 76 176 84 184
rect 252 396 260 404
rect 220 316 228 324
rect 380 696 388 704
rect 460 696 468 704
rect 492 696 500 704
rect 638 806 646 814
rect 652 806 660 814
rect 666 806 674 814
rect 748 736 756 744
rect 540 716 548 724
rect 700 716 708 724
rect 556 696 564 704
rect 476 676 484 684
rect 460 636 468 644
rect 364 596 372 604
rect 428 616 436 624
rect 348 576 356 584
rect 412 576 420 584
rect 364 556 372 564
rect 508 676 516 684
rect 572 676 580 684
rect 540 656 548 664
rect 732 676 740 684
rect 588 656 596 664
rect 668 656 676 664
rect 556 636 564 644
rect 748 636 756 644
rect 524 556 532 564
rect 380 536 388 544
rect 508 516 516 524
rect 572 516 580 524
rect 700 516 708 524
rect 604 476 612 484
rect 348 396 356 404
rect 638 406 646 414
rect 652 406 660 414
rect 666 406 674 414
rect 556 336 564 344
rect 716 336 724 344
rect 556 316 564 324
rect 140 136 148 144
rect 268 136 276 144
rect 524 276 532 284
rect 636 296 644 304
rect 924 996 932 1004
rect 988 976 996 984
rect 860 956 868 964
rect 892 936 900 944
rect 1116 1316 1124 1324
rect 1212 1236 1220 1244
rect 1260 1236 1268 1244
rect 1372 1696 1380 1704
rect 1484 1896 1492 1904
rect 1516 1896 1524 1904
rect 1468 1776 1476 1784
rect 1404 1516 1412 1524
rect 1404 1496 1412 1504
rect 1356 1476 1364 1484
rect 1468 1496 1476 1504
rect 1452 1476 1460 1484
rect 1468 1476 1476 1484
rect 1436 1236 1444 1244
rect 1244 1176 1252 1184
rect 1436 1176 1444 1184
rect 1084 976 1092 984
rect 1068 936 1076 944
rect 1100 956 1108 964
rect 1132 936 1140 944
rect 1212 916 1220 924
rect 1308 1156 1316 1164
rect 1468 1156 1476 1164
rect 1324 1136 1332 1144
rect 1500 1856 1508 1864
rect 1532 1856 1540 1864
rect 1516 1836 1524 1844
rect 1550 1806 1558 1814
rect 1564 1806 1572 1814
rect 1578 1806 1586 1814
rect 1580 1756 1588 1764
rect 1596 1716 1604 1724
rect 1516 1696 1524 1704
rect 1612 1496 1620 1504
rect 1500 1476 1508 1484
rect 1612 1476 1620 1484
rect 1820 1996 1828 2004
rect 1868 1996 1876 2004
rect 1676 1836 1684 1844
rect 1676 1796 1684 1804
rect 1772 1796 1780 1804
rect 1644 1776 1652 1784
rect 1740 1756 1748 1764
rect 1660 1716 1668 1724
rect 1836 1756 1844 1764
rect 2044 1896 2052 1904
rect 2140 1896 2148 1904
rect 2188 1896 2196 1904
rect 2236 1896 2244 1904
rect 2092 1876 2100 1884
rect 2156 1856 2164 1864
rect 2076 1756 2084 1764
rect 1884 1716 1892 1724
rect 1948 1716 1956 1724
rect 1756 1496 1764 1504
rect 1804 1496 1812 1504
rect 1980 1496 1988 1504
rect 1550 1406 1558 1414
rect 1564 1406 1572 1414
rect 1578 1406 1586 1414
rect 1772 1476 1780 1484
rect 1804 1476 1812 1484
rect 1836 1456 1844 1464
rect 1804 1436 1812 1444
rect 1836 1436 1844 1444
rect 1676 1396 1684 1404
rect 1740 1396 1748 1404
rect 1500 1336 1508 1344
rect 1644 1336 1652 1344
rect 2012 1396 2020 1404
rect 1580 1316 1588 1324
rect 1900 1316 1908 1324
rect 1644 1176 1652 1184
rect 1484 1136 1492 1144
rect 1500 1136 1508 1144
rect 1404 1116 1412 1124
rect 1452 1116 1460 1124
rect 1276 1096 1284 1104
rect 1388 1096 1396 1104
rect 1420 1096 1428 1104
rect 1260 916 1268 924
rect 1164 896 1172 904
rect 1500 1096 1508 1104
rect 1564 1096 1572 1104
rect 1324 1056 1332 1064
rect 1532 1056 1540 1064
rect 1356 1036 1364 1044
rect 1356 996 1364 1004
rect 1308 916 1316 924
rect 1180 816 1188 824
rect 1084 796 1092 804
rect 1180 796 1188 804
rect 780 696 788 704
rect 1132 696 1134 704
rect 1134 696 1140 704
rect 796 656 804 664
rect 796 336 804 344
rect 748 316 756 324
rect 764 316 772 324
rect 796 316 804 324
rect 940 676 948 684
rect 1212 676 1220 684
rect 972 636 980 644
rect 1036 616 1044 624
rect 876 596 884 604
rect 1020 556 1028 564
rect 1004 536 1012 544
rect 1100 536 1108 544
rect 1068 496 1076 504
rect 908 476 916 484
rect 844 336 852 344
rect 828 296 836 304
rect 1004 416 1012 424
rect 1004 356 1012 364
rect 924 336 932 344
rect 1052 356 1060 364
rect 1084 356 1092 364
rect 1116 516 1124 524
rect 1132 496 1140 504
rect 1148 476 1156 484
rect 1212 516 1220 524
rect 1836 1156 1844 1164
rect 1740 1116 1748 1124
rect 1948 1216 1956 1224
rect 1996 1216 2004 1224
rect 1916 1136 1924 1144
rect 1868 1116 1876 1124
rect 1900 1116 1908 1124
rect 1708 1096 1716 1104
rect 1820 1096 1828 1104
rect 1852 1096 1860 1104
rect 1980 1096 1988 1104
rect 2092 1096 2100 1104
rect 1692 1076 1700 1084
rect 1676 1056 1684 1064
rect 1564 1036 1572 1044
rect 1660 1036 1668 1044
rect 1550 1006 1558 1014
rect 1564 1006 1572 1014
rect 1578 1006 1586 1014
rect 1452 996 1460 1004
rect 1516 956 1524 964
rect 1388 916 1396 924
rect 1436 896 1444 904
rect 1548 936 1556 944
rect 1612 916 1620 924
rect 1260 676 1268 684
rect 1292 676 1300 684
rect 1244 616 1252 624
rect 1276 516 1284 524
rect 1196 496 1204 504
rect 1212 496 1220 504
rect 1164 356 1172 364
rect 1132 336 1140 344
rect 1164 336 1172 344
rect 812 276 820 284
rect 956 276 964 284
rect 892 256 900 264
rect 540 136 548 144
rect 988 296 996 304
rect 1020 296 1028 304
rect 972 256 980 264
rect 1116 316 1124 324
rect 1212 456 1220 464
rect 1228 416 1236 424
rect 1100 276 1108 284
rect 1116 276 1124 284
rect 1100 256 1108 264
rect 1180 256 1188 264
rect 1196 256 1204 264
rect 1260 176 1268 184
rect 1420 636 1428 644
rect 1420 536 1428 544
rect 1452 536 1460 544
rect 1340 476 1348 484
rect 1308 176 1316 184
rect 1260 156 1268 164
rect 1292 156 1300 164
rect 908 136 916 144
rect 1612 676 1620 684
rect 1532 636 1540 644
rect 1644 636 1652 644
rect 1550 606 1558 614
rect 1564 606 1572 614
rect 1578 606 1586 614
rect 1644 576 1652 584
rect 1676 536 1684 544
rect 1708 536 1716 544
rect 1756 1036 1764 1044
rect 1852 1056 1860 1064
rect 1964 1036 1972 1044
rect 1804 1016 1812 1024
rect 1900 956 1908 964
rect 1772 936 1780 944
rect 1772 916 1780 924
rect 1868 836 1876 844
rect 1916 836 1924 844
rect 1884 756 1892 764
rect 1948 736 1956 744
rect 2044 1056 2052 1064
rect 2108 1056 2116 1064
rect 2124 1036 2132 1044
rect 2028 956 2036 964
rect 2092 1016 2100 1024
rect 2140 956 2148 964
rect 2172 1456 2180 1464
rect 2188 1076 2196 1084
rect 2188 1056 2196 1064
rect 2172 956 2180 964
rect 2156 936 2164 944
rect 2076 916 2084 924
rect 2060 796 2068 804
rect 2060 736 2068 744
rect 1852 716 1860 724
rect 1900 716 1908 724
rect 1980 716 1988 724
rect 1756 696 1764 704
rect 1852 696 1860 704
rect 2092 896 2100 904
rect 2156 916 2164 924
rect 2172 916 2180 924
rect 2156 896 2164 904
rect 2124 876 2132 884
rect 2252 1856 2260 1864
rect 2252 1496 2260 1504
rect 2252 1136 2260 1144
rect 2220 1096 2228 1104
rect 2204 936 2212 944
rect 2220 916 2228 924
rect 2172 816 2180 824
rect 2108 756 2116 764
rect 2124 736 2132 744
rect 2172 736 2180 744
rect 2092 716 2100 724
rect 1980 696 1988 704
rect 2028 696 2036 704
rect 2076 696 2084 704
rect 2108 696 2116 704
rect 2124 696 2132 704
rect 2172 696 2180 704
rect 1836 676 1844 684
rect 1900 676 1908 684
rect 1852 656 1860 664
rect 1804 636 1812 644
rect 1772 536 1780 544
rect 1836 536 1844 544
rect 1660 516 1668 524
rect 1772 516 1780 524
rect 1820 516 1828 524
rect 1804 476 1812 484
rect 1724 456 1732 464
rect 1692 436 1700 444
rect 1420 236 1428 244
rect 1356 176 1364 184
rect 1372 176 1380 184
rect 1468 176 1476 184
rect 1452 156 1460 164
rect 1404 136 1412 144
rect 1468 136 1476 144
rect 1612 276 1620 284
rect 1676 276 1684 284
rect 1550 206 1558 214
rect 1564 206 1572 214
rect 1578 206 1586 214
rect 1628 256 1636 264
rect 1692 256 1700 264
rect 1708 256 1716 264
rect 1612 196 1620 204
rect 1564 176 1572 184
rect 1532 156 1540 164
rect 1756 276 1764 284
rect 1772 276 1780 284
rect 1804 276 1812 284
rect 1772 256 1780 264
rect 1836 496 1844 504
rect 1868 636 1876 644
rect 1996 676 2004 684
rect 2076 676 2084 684
rect 2156 676 2164 684
rect 1964 656 1972 664
rect 2012 656 2020 664
rect 2028 656 2036 664
rect 2060 656 2068 664
rect 2124 656 2132 664
rect 1900 576 1908 584
rect 1996 576 2004 584
rect 1980 536 1988 544
rect 1868 516 1876 524
rect 1884 476 1892 484
rect 1820 216 1828 224
rect 2156 636 2164 644
rect 2140 576 2148 584
rect 2108 556 2116 564
rect 2044 536 2052 544
rect 2044 516 2052 524
rect 2108 496 2116 504
rect 1900 356 1908 364
rect 1948 356 1956 364
rect 1932 336 1940 344
rect 1948 336 1956 344
rect 1916 316 1924 324
rect 1980 316 1988 324
rect 2108 436 2116 444
rect 2012 296 2020 304
rect 2060 296 2068 304
rect 2108 296 2116 304
rect 1884 256 1892 264
rect 2028 276 2036 284
rect 1996 256 2004 264
rect 1868 236 1876 244
rect 1932 236 1940 244
rect 1852 196 1860 204
rect 1724 136 1732 144
rect 2044 256 2052 264
rect 2092 236 2100 244
rect 2108 176 2116 184
rect 2140 536 2148 544
rect 2220 876 2228 884
rect 2204 856 2212 864
rect 2236 816 2244 824
rect 2204 716 2212 724
rect 2220 576 2228 584
rect 2172 556 2180 564
rect 2188 536 2196 544
rect 2252 676 2260 684
rect 2156 336 2164 344
rect 2252 336 2260 344
rect 2172 296 2180 304
rect 2156 256 2164 264
rect 2204 256 2212 264
rect 2204 216 2212 224
rect 2060 156 2068 164
rect 2188 156 2196 164
rect 364 116 372 124
rect 444 116 452 124
rect 1212 116 1220 124
rect 1340 116 1348 124
rect 1356 116 1364 124
rect 1420 116 1428 124
rect 1516 116 1524 124
rect 1788 116 1796 124
rect 12 96 20 104
rect 1516 96 1524 104
rect 1612 96 1620 104
rect 2092 96 2100 104
rect 2124 96 2132 104
rect 2252 96 2260 104
rect 812 16 820 24
rect 844 16 852 24
rect 638 6 646 14
rect 652 6 660 14
rect 666 6 674 14
<< metal3 >>
rect 632 2014 680 2016
rect 632 2006 636 2014
rect 646 2006 652 2014
rect 660 2006 666 2014
rect 676 2006 680 2014
rect 632 2004 680 2006
rect 1828 1997 1868 2003
rect 1460 1917 1500 1923
rect -19 1897 12 1903
rect 900 1897 1004 1903
rect 1492 1897 1516 1903
rect 2052 1897 2099 1903
rect 2093 1884 2099 1897
rect 2148 1897 2188 1903
rect 2196 1897 2236 1903
rect 148 1877 268 1883
rect 916 1877 1132 1883
rect 1524 1877 2092 1883
rect 1508 1857 1532 1863
rect 2164 1857 2252 1863
rect 2260 1857 2291 1863
rect 532 1837 572 1843
rect 1524 1837 1676 1843
rect 180 1817 732 1823
rect 740 1817 812 1823
rect 820 1817 1052 1823
rect 1060 1817 1100 1823
rect 1108 1817 1340 1823
rect 1348 1817 1516 1823
rect 1544 1814 1592 1816
rect 1544 1806 1548 1814
rect 1558 1806 1564 1814
rect 1572 1806 1578 1814
rect 1588 1806 1592 1814
rect 1544 1804 1592 1806
rect 372 1797 492 1803
rect 500 1797 812 1803
rect 820 1797 972 1803
rect 1060 1797 1308 1803
rect 1684 1797 1772 1803
rect 404 1777 780 1783
rect 1284 1777 1308 1783
rect 1428 1777 1468 1783
rect 1476 1777 1644 1783
rect 244 1757 364 1763
rect 372 1757 684 1763
rect 804 1757 844 1763
rect 1444 1757 1580 1763
rect 1748 1757 1836 1763
rect 1844 1757 2076 1763
rect 717 1737 764 1743
rect 717 1724 723 1737
rect 820 1737 908 1743
rect 580 1717 716 1723
rect 756 1717 828 1723
rect 1188 1717 1228 1723
rect 1284 1717 1340 1723
rect 1364 1717 1388 1723
rect 1604 1717 1660 1723
rect 1892 1717 1948 1723
rect -19 1697 12 1703
rect 1172 1697 1260 1703
rect 1268 1697 1372 1703
rect 1380 1697 1516 1703
rect 612 1677 1292 1683
rect 52 1657 204 1663
rect 212 1657 540 1663
rect 1060 1617 1132 1623
rect 632 1614 680 1616
rect 632 1606 636 1614
rect 646 1606 652 1614
rect 660 1606 666 1614
rect 676 1606 680 1614
rect 632 1604 680 1606
rect 1332 1517 1404 1523
rect -19 1497 12 1503
rect 372 1497 396 1503
rect 452 1497 524 1503
rect 532 1497 748 1503
rect 868 1497 972 1503
rect 1300 1497 1404 1503
rect 1412 1497 1468 1503
rect 1620 1497 1756 1503
rect 1812 1497 1980 1503
rect 2260 1497 2291 1503
rect 148 1477 268 1483
rect 404 1477 412 1483
rect 468 1477 540 1483
rect 1108 1477 1308 1483
rect 1364 1477 1452 1483
rect 1476 1477 1500 1483
rect 1524 1477 1612 1483
rect 1780 1477 1804 1483
rect 244 1457 364 1463
rect 436 1457 476 1463
rect 964 1457 1100 1463
rect 1108 1457 1132 1463
rect 1140 1457 1244 1463
rect 1844 1457 2172 1463
rect 1812 1437 1836 1443
rect 756 1417 844 1423
rect 1544 1414 1592 1416
rect 1544 1406 1548 1414
rect 1558 1406 1564 1414
rect 1572 1406 1578 1414
rect 1588 1406 1592 1414
rect 1544 1404 1592 1406
rect 1684 1397 1740 1403
rect 1748 1397 2012 1403
rect 52 1377 204 1383
rect 212 1377 540 1383
rect 596 1357 748 1363
rect 404 1337 492 1343
rect 756 1337 796 1343
rect 1508 1337 1644 1343
rect 532 1317 556 1323
rect 564 1317 604 1323
rect 788 1317 828 1323
rect 1012 1317 1116 1323
rect 1588 1317 1900 1323
rect -19 1297 12 1303
rect 932 1297 1068 1303
rect 1076 1297 1516 1303
rect 292 1277 396 1283
rect 404 1277 588 1283
rect 596 1277 876 1283
rect 372 1237 540 1243
rect 1220 1237 1260 1243
rect 1268 1237 1436 1243
rect 132 1217 156 1223
rect 164 1217 316 1223
rect 1956 1217 1996 1223
rect 632 1214 680 1216
rect 632 1206 636 1214
rect 646 1206 652 1214
rect 660 1206 666 1214
rect 676 1206 680 1214
rect 632 1204 680 1206
rect 1252 1177 1436 1183
rect 1444 1177 1644 1183
rect 1316 1157 1468 1163
rect 1476 1157 1804 1163
rect 1812 1157 1836 1163
rect -19 1137 12 1143
rect 804 1137 1324 1143
rect 1332 1137 1484 1143
rect 1508 1137 1916 1143
rect 2260 1137 2291 1143
rect 180 1117 252 1123
rect 797 1123 803 1136
rect 260 1117 803 1123
rect 1412 1117 1443 1123
rect -19 1097 60 1103
rect 372 1097 572 1103
rect 676 1097 988 1103
rect 1284 1097 1388 1103
rect 1396 1097 1420 1103
rect 1437 1103 1443 1117
rect 1460 1117 1740 1123
rect 1748 1117 1868 1123
rect 1908 1117 2291 1123
rect 1437 1097 1500 1103
rect 1572 1097 1708 1103
rect 1828 1097 1852 1103
rect 1860 1097 1980 1103
rect 2100 1097 2220 1103
rect 2285 1097 2291 1117
rect 116 1077 220 1083
rect 228 1077 380 1083
rect 1533 1077 1692 1083
rect 1533 1064 1539 1077
rect 1700 1077 2188 1083
rect 52 1057 140 1063
rect 228 1057 268 1063
rect 308 1057 444 1063
rect 548 1057 764 1063
rect 772 1057 796 1063
rect 1332 1057 1532 1063
rect 1684 1057 1852 1063
rect 2052 1057 2108 1063
rect 2116 1057 2188 1063
rect 356 1037 412 1043
rect 1364 1037 1564 1043
rect 1668 1037 1756 1043
rect 1972 1037 2124 1043
rect 788 1017 908 1023
rect 1812 1017 2092 1023
rect 1544 1014 1592 1016
rect 1544 1006 1548 1014
rect 1558 1006 1564 1014
rect 1572 1006 1578 1014
rect 1588 1006 1592 1014
rect 1544 1004 1592 1006
rect 884 997 924 1003
rect 1364 997 1452 1003
rect 388 977 476 983
rect 996 977 1084 983
rect 404 957 467 963
rect 461 944 467 957
rect 868 957 1100 963
rect 1524 957 1900 963
rect 2036 957 2140 963
rect 2148 957 2172 963
rect 2180 957 2252 963
rect 292 937 412 943
rect 468 937 572 943
rect 580 937 700 943
rect 756 937 892 943
rect 1076 937 1132 943
rect 1140 937 1164 943
rect 1556 937 1772 943
rect 2196 937 2204 943
rect 452 917 460 923
rect 468 917 588 923
rect 1220 917 1260 923
rect 1268 917 1308 923
rect 1316 917 1388 923
rect 1620 917 1772 923
rect 2084 917 2156 923
rect 2180 917 2220 923
rect -19 897 364 903
rect 1172 897 1436 903
rect 2100 897 2156 903
rect 2036 877 2124 883
rect 2132 877 2220 883
rect 2212 857 2220 863
rect 1876 837 1916 843
rect 1044 817 1180 823
rect 2180 817 2236 823
rect 632 814 680 816
rect 632 806 636 814
rect 646 806 652 814
rect 660 806 666 814
rect 676 806 680 814
rect 632 804 680 806
rect 1092 797 1180 803
rect 1892 757 2108 763
rect 436 737 748 743
rect 1956 737 2060 743
rect 2132 737 2172 743
rect 548 717 700 723
rect 1652 717 1852 723
rect 1908 717 1980 723
rect 1988 717 2092 723
rect 2212 717 2291 723
rect 388 697 460 703
rect 500 697 556 703
rect 788 697 1132 703
rect 1764 697 1852 703
rect 1988 697 2028 703
rect 2084 697 2108 703
rect 2132 697 2172 703
rect 36 677 476 683
rect 516 677 572 683
rect 740 677 940 683
rect 1220 677 1260 683
rect 1268 677 1292 683
rect 1620 677 1644 683
rect 1844 677 1900 683
rect 2004 677 2076 683
rect 2084 677 2156 683
rect 2164 677 2252 683
rect 2260 677 2291 683
rect 548 657 588 663
rect 676 657 796 663
rect 1812 657 1852 663
rect 1860 657 1964 663
rect 2020 657 2028 663
rect 2036 657 2060 663
rect 2068 657 2124 663
rect 468 637 556 643
rect 756 637 972 643
rect 1428 637 1532 643
rect 1540 637 1644 643
rect 1812 637 1868 643
rect 2164 637 2188 643
rect 228 617 268 623
rect 292 617 428 623
rect 1044 617 1244 623
rect 1544 614 1592 616
rect 1544 606 1548 614
rect 1558 606 1564 614
rect 1572 606 1578 614
rect 1588 606 1592 614
rect 1544 604 1592 606
rect 228 597 364 603
rect 196 577 236 583
rect 356 577 412 583
rect 1652 577 1900 583
rect 1908 577 1996 583
rect 2148 577 2220 583
rect 2228 577 2291 583
rect 52 557 220 563
rect 324 557 364 563
rect 372 557 524 563
rect 1028 557 1036 563
rect 2116 557 2172 563
rect -19 537 12 543
rect 100 537 380 543
rect 1012 537 1100 543
rect 1108 537 1420 543
rect 1460 537 1676 543
rect 1716 537 1772 543
rect 1844 537 1980 543
rect 2052 537 2140 543
rect 2196 537 2291 543
rect 36 517 124 523
rect 180 517 188 523
rect 196 517 508 523
rect 580 517 700 523
rect 1124 517 1212 523
rect 1284 517 1660 523
rect 1780 517 1820 523
rect 1828 517 1868 523
rect 1981 523 1987 536
rect 1981 517 2044 523
rect 2052 517 2060 523
rect -19 497 60 503
rect 180 497 204 503
rect 1076 497 1132 503
rect 1140 497 1196 503
rect 1220 497 1836 503
rect 2116 497 2291 503
rect 244 477 300 483
rect 308 477 604 483
rect 612 477 908 483
rect 1156 477 1340 483
rect 1812 477 1884 483
rect 1220 457 1724 463
rect 1700 437 2108 443
rect 1012 417 1228 423
rect 632 414 680 416
rect 632 406 636 414
rect 646 406 652 414
rect 660 406 666 414
rect 676 406 680 414
rect 632 404 680 406
rect 260 397 348 403
rect 68 377 92 383
rect 845 357 1004 363
rect 845 344 851 357
rect 1060 357 1084 363
rect 1092 357 1164 363
rect 1908 357 1948 363
rect 724 337 796 343
rect 804 337 844 343
rect 932 337 1132 343
rect 1172 337 1932 343
rect 1956 337 2156 343
rect 2228 337 2252 343
rect 2260 337 2291 343
rect 228 317 236 323
rect 244 317 556 323
rect 564 317 748 323
rect 772 317 796 323
rect 804 317 1116 323
rect 1924 317 1980 323
rect 644 297 828 303
rect 996 297 1020 303
rect 2020 297 2028 303
rect 2036 297 2060 303
rect 2116 297 2172 303
rect 2196 297 2291 303
rect 532 277 812 283
rect 964 277 1100 283
rect 1124 277 1612 283
rect 1684 277 1756 283
rect 1780 277 1804 283
rect 2036 277 2156 283
rect 900 257 972 263
rect 1108 257 1180 263
rect 1204 257 1628 263
rect 1636 257 1692 263
rect 1716 257 1772 263
rect 1780 257 1884 263
rect 2004 257 2044 263
rect 2164 257 2188 263
rect 2212 257 2252 263
rect 2260 257 2291 263
rect 1428 237 1868 243
rect 1940 237 2092 243
rect 1828 217 2204 223
rect 1544 214 1592 216
rect 1544 206 1548 214
rect 1558 206 1564 214
rect 1572 206 1578 214
rect 1588 206 1592 214
rect 1544 204 1592 206
rect 1620 197 1852 203
rect 20 177 76 183
rect 1268 177 1308 183
rect 1316 177 1356 183
rect 1380 177 1468 183
rect 1572 177 2108 183
rect 1268 157 1292 163
rect 1460 157 1532 163
rect 2068 157 2188 163
rect 148 137 268 143
rect 548 137 556 143
rect 916 137 1404 143
rect 1476 137 1724 143
rect 372 117 444 123
rect 1220 117 1340 123
rect 1364 117 1420 123
rect 1524 117 1788 123
rect -19 97 12 103
rect 1524 97 1612 103
rect 2100 97 2124 103
rect 2260 97 2291 103
rect 820 17 844 23
rect 632 14 680 16
rect 632 6 636 14
rect 646 6 652 14
rect 660 6 666 14
rect 676 6 680 14
rect 632 4 680 6
<< m4contact >>
rect 636 2006 638 2014
rect 638 2006 644 2014
rect 652 2006 660 2014
rect 668 2006 674 2014
rect 674 2006 676 2014
rect 1516 1876 1524 1884
rect 812 1816 820 1824
rect 1516 1816 1524 1824
rect 1548 1806 1550 1814
rect 1550 1806 1556 1814
rect 1564 1806 1572 1814
rect 1580 1806 1586 1814
rect 1586 1806 1588 1814
rect 1164 1696 1172 1704
rect 636 1606 638 1614
rect 638 1606 644 1614
rect 652 1606 660 1614
rect 668 1606 674 1614
rect 674 1606 676 1614
rect 172 1596 180 1604
rect 396 1476 404 1484
rect 1516 1476 1524 1484
rect 1548 1406 1550 1414
rect 1550 1406 1556 1414
rect 1564 1406 1572 1414
rect 1580 1406 1586 1414
rect 1586 1406 1588 1414
rect 812 1336 820 1344
rect 172 1316 180 1324
rect 1516 1296 1524 1304
rect 396 1276 404 1284
rect 636 1206 638 1214
rect 638 1206 644 1214
rect 652 1206 660 1214
rect 668 1206 674 1214
rect 674 1206 676 1214
rect 1804 1156 1812 1164
rect 1548 1006 1550 1014
rect 1550 1006 1556 1014
rect 1564 1006 1572 1014
rect 1580 1006 1586 1014
rect 1586 1006 1588 1014
rect 876 996 884 1004
rect 2252 956 2260 964
rect 1164 936 1172 944
rect 2156 936 2164 944
rect 2188 936 2196 944
rect 2028 876 2036 884
rect 2220 856 2228 864
rect 1036 816 1044 824
rect 636 806 638 814
rect 638 806 644 814
rect 652 806 660 814
rect 668 806 674 814
rect 674 806 676 814
rect 2060 796 2068 804
rect 1644 716 1652 724
rect 1644 676 1652 684
rect 1804 656 1812 664
rect 2188 636 2196 644
rect 1548 606 1550 614
rect 1550 606 1556 614
rect 1564 606 1572 614
rect 1580 606 1586 614
rect 1586 606 1588 614
rect 876 596 884 604
rect 236 576 244 584
rect 1036 556 1044 564
rect 172 516 180 524
rect 2060 516 2068 524
rect 636 406 638 414
rect 638 406 644 414
rect 652 406 660 414
rect 668 406 674 414
rect 674 406 676 414
rect 556 336 564 344
rect 2220 336 2228 344
rect 236 316 244 324
rect 2028 296 2036 304
rect 2188 296 2196 304
rect 2156 276 2164 284
rect 2188 256 2196 264
rect 2252 256 2260 264
rect 1548 206 1550 214
rect 1550 206 1556 214
rect 1564 206 1572 214
rect 1580 206 1586 214
rect 1586 206 1588 214
rect 556 136 564 144
rect 636 6 638 14
rect 638 6 644 14
rect 652 6 660 14
rect 668 6 674 14
rect 674 6 676 14
<< metal4 >>
rect 632 2014 680 2040
rect 632 2006 636 2014
rect 644 2006 652 2014
rect 660 2006 668 2014
rect 676 2006 680 2014
rect 632 1614 680 2006
rect 1514 1884 1526 1886
rect 1514 1876 1516 1884
rect 1524 1876 1526 1884
rect 632 1606 636 1614
rect 644 1606 652 1614
rect 660 1606 668 1614
rect 676 1606 680 1614
rect 170 1604 182 1606
rect 170 1596 172 1604
rect 180 1596 182 1604
rect 170 1324 182 1596
rect 170 1316 172 1324
rect 180 1316 182 1324
rect 170 524 182 1316
rect 394 1484 406 1486
rect 394 1476 396 1484
rect 404 1476 406 1484
rect 394 1284 406 1476
rect 394 1276 396 1284
rect 404 1276 406 1284
rect 394 1274 406 1276
rect 632 1214 680 1606
rect 810 1824 822 1826
rect 810 1816 812 1824
rect 820 1816 822 1824
rect 810 1344 822 1816
rect 1514 1824 1526 1876
rect 1514 1816 1516 1824
rect 1524 1816 1526 1824
rect 1514 1814 1526 1816
rect 1544 1814 1592 2040
rect 1544 1806 1548 1814
rect 1556 1806 1564 1814
rect 1572 1806 1580 1814
rect 1588 1806 1592 1814
rect 810 1336 812 1344
rect 820 1336 822 1344
rect 810 1334 822 1336
rect 1162 1704 1174 1706
rect 1162 1696 1164 1704
rect 1172 1696 1174 1704
rect 632 1206 636 1214
rect 644 1206 652 1214
rect 660 1206 668 1214
rect 676 1206 680 1214
rect 632 814 680 1206
rect 632 806 636 814
rect 644 806 652 814
rect 660 806 668 814
rect 676 806 680 814
rect 170 516 172 524
rect 180 516 182 524
rect 170 514 182 516
rect 234 584 246 586
rect 234 576 236 584
rect 244 576 246 584
rect 234 324 246 576
rect 632 414 680 806
rect 874 1004 886 1006
rect 874 996 876 1004
rect 884 996 886 1004
rect 874 604 886 996
rect 1162 944 1174 1696
rect 1514 1484 1526 1486
rect 1514 1476 1516 1484
rect 1524 1476 1526 1484
rect 1514 1304 1526 1476
rect 1514 1296 1516 1304
rect 1524 1296 1526 1304
rect 1514 1294 1526 1296
rect 1544 1414 1592 1806
rect 1544 1406 1548 1414
rect 1556 1406 1564 1414
rect 1572 1406 1580 1414
rect 1588 1406 1592 1414
rect 1162 936 1164 944
rect 1172 936 1174 944
rect 1162 934 1174 936
rect 1544 1014 1592 1406
rect 1544 1006 1548 1014
rect 1556 1006 1564 1014
rect 1572 1006 1580 1014
rect 1588 1006 1592 1014
rect 874 596 876 604
rect 884 596 886 604
rect 874 594 886 596
rect 1034 824 1046 826
rect 1034 816 1036 824
rect 1044 816 1046 824
rect 1034 564 1046 816
rect 1034 556 1036 564
rect 1044 556 1046 564
rect 1034 554 1046 556
rect 1544 614 1592 1006
rect 1802 1164 1814 1166
rect 1802 1156 1804 1164
rect 1812 1156 1814 1164
rect 1642 724 1654 726
rect 1642 716 1644 724
rect 1652 716 1654 724
rect 1642 684 1654 716
rect 1642 676 1644 684
rect 1652 676 1654 684
rect 1642 674 1654 676
rect 1802 664 1814 1156
rect 2250 964 2262 966
rect 2250 956 2252 964
rect 2260 956 2262 964
rect 2154 944 2166 946
rect 2154 936 2156 944
rect 2164 936 2166 944
rect 1802 656 1804 664
rect 1812 656 1814 664
rect 1802 654 1814 656
rect 2026 884 2038 886
rect 2026 876 2028 884
rect 2036 876 2038 884
rect 1544 606 1548 614
rect 1556 606 1564 614
rect 1572 606 1580 614
rect 1588 606 1592 614
rect 632 406 636 414
rect 644 406 652 414
rect 660 406 668 414
rect 676 406 680 414
rect 234 316 236 324
rect 244 316 246 324
rect 234 314 246 316
rect 554 344 566 346
rect 554 336 556 344
rect 564 336 566 344
rect 554 144 566 336
rect 554 136 556 144
rect 564 136 566 144
rect 554 134 566 136
rect 632 14 680 406
rect 632 6 636 14
rect 644 6 652 14
rect 660 6 668 14
rect 676 6 680 14
rect 632 -40 680 6
rect 1544 214 1592 606
rect 2026 304 2038 876
rect 2058 804 2070 806
rect 2058 796 2060 804
rect 2068 796 2070 804
rect 2058 524 2070 796
rect 2058 516 2060 524
rect 2068 516 2070 524
rect 2058 514 2070 516
rect 2026 296 2028 304
rect 2036 296 2038 304
rect 2026 294 2038 296
rect 2154 284 2166 936
rect 2186 944 2198 946
rect 2186 936 2188 944
rect 2196 936 2198 944
rect 2186 644 2198 936
rect 2186 636 2188 644
rect 2196 636 2198 644
rect 2186 634 2198 636
rect 2218 864 2230 866
rect 2218 856 2220 864
rect 2228 856 2230 864
rect 2218 344 2230 856
rect 2218 336 2220 344
rect 2228 336 2230 344
rect 2218 334 2230 336
rect 2154 276 2156 284
rect 2164 276 2166 284
rect 2154 274 2166 276
rect 2186 304 2198 306
rect 2186 296 2188 304
rect 2196 296 2198 304
rect 2186 264 2198 296
rect 2186 256 2188 264
rect 2196 256 2198 264
rect 2186 254 2198 256
rect 2250 264 2262 956
rect 2250 256 2252 264
rect 2260 256 2262 264
rect 2250 254 2262 256
rect 1544 206 1548 214
rect 1556 206 1564 214
rect 1572 206 1580 214
rect 1588 206 1592 214
rect 1544 -40 1592 206
use BUFX2  BUFX2_25
timestamp 1560284232
transform -1 0 56 0 1 1810
box 0 0 48 200
use DFFSR  DFFSR_30
timestamp 1560284232
transform -1 0 408 0 1 1810
box 0 0 352 200
use BUFX2  BUFX2_21
timestamp 1560284232
transform -1 0 456 0 1 1810
box 0 0 48 200
use FILL  FILL_9_0_0
timestamp 1560284232
transform -1 0 472 0 1 1810
box 0 0 16 200
use FILL  FILL_9_0_1
timestamp 1560284232
transform -1 0 488 0 1 1810
box 0 0 16 200
use FILL  FILL_9_0_2
timestamp 1560284232
transform -1 0 504 0 1 1810
box 0 0 16 200
use DFFSR  DFFSR_26
timestamp 1560284232
transform -1 0 856 0 1 1810
box 0 0 352 200
use BUFX2  BUFX2_20
timestamp 1560284232
transform -1 0 904 0 1 1810
box 0 0 48 200
use BUFX2  BUFX2_28
timestamp 1560284232
transform 1 0 904 0 1 1810
box 0 0 48 200
use BUFX2  BUFX2_23
timestamp 1560284232
transform 1 0 952 0 1 1810
box 0 0 48 200
use INVX1  INVX1_5
timestamp 1560284232
transform 1 0 1000 0 1 1810
box 0 0 32 200
use AOI21X1  AOI21X1_1
timestamp 1560284232
transform 1 0 1032 0 1 1810
box 0 0 64 200
use NOR2X1  NOR2X1_4
timestamp 1560284232
transform -1 0 1144 0 1 1810
box 0 0 48 200
use DFFSR  DFFSR_27
timestamp 1560284232
transform 1 0 1144 0 1 1810
box 0 0 352 200
use NAND3X1  NAND3X1_3
timestamp 1560284232
transform 1 0 1496 0 1 1810
box 0 0 64 200
use FILL  FILL_9_1_0
timestamp 1560284232
transform -1 0 1576 0 1 1810
box 0 0 16 200
use FILL  FILL_9_1_1
timestamp 1560284232
transform -1 0 1592 0 1 1810
box 0 0 16 200
use FILL  FILL_9_1_2
timestamp 1560284232
transform -1 0 1608 0 1 1810
box 0 0 16 200
use BUFX2  BUFX2_22
timestamp 1560284232
transform -1 0 1656 0 1 1810
box 0 0 48 200
use DFFSR  DFFSR_6
timestamp 1560284232
transform -1 0 2008 0 1 1810
box 0 0 352 200
use NOR2X1  NOR2X1_5
timestamp 1560284232
transform 1 0 2008 0 1 1810
box 0 0 48 200
use AOI21X1  AOI21X1_2
timestamp 1560284232
transform -1 0 2120 0 1 1810
box 0 0 64 200
use INVX1  INVX1_21
timestamp 1560284232
transform -1 0 2152 0 1 1810
box 0 0 32 200
use BUFX2  BUFX2_19
timestamp 1560284232
transform -1 0 2200 0 1 1810
box 0 0 48 200
use INVX1  INVX1_32
timestamp 1560284232
transform -1 0 2232 0 1 1810
box 0 0 32 200
use FILL  FILL_10_1
timestamp 1560284232
transform 1 0 2232 0 1 1810
box 0 0 16 200
use FILL  FILL_10_2
timestamp 1560284232
transform 1 0 2248 0 1 1810
box 0 0 16 200
use BUFX2  BUFX2_29
timestamp 1560284232
transform -1 0 56 0 -1 1810
box 0 0 48 200
use INVX1  INVX1_15
timestamp 1560284232
transform 1 0 56 0 -1 1810
box 0 0 32 200
use MUX2X1  MUX2X1_5
timestamp 1560284232
transform -1 0 184 0 -1 1810
box 0 0 96 200
use DFFSR  DFFSR_17
timestamp 1560284232
transform -1 0 536 0 -1 1810
box 0 0 352 200
use INVX1  INVX1_8
timestamp 1560284232
transform 1 0 536 0 -1 1810
box 0 0 32 200
use INVX1  INVX1_7
timestamp 1560284232
transform 1 0 568 0 -1 1810
box 0 0 32 200
use FILL  FILL_8_0_0
timestamp 1560284232
transform -1 0 616 0 -1 1810
box 0 0 16 200
use FILL  FILL_8_0_1
timestamp 1560284232
transform -1 0 632 0 -1 1810
box 0 0 16 200
use FILL  FILL_8_0_2
timestamp 1560284232
transform -1 0 648 0 -1 1810
box 0 0 16 200
use MUX2X1  MUX2X1_1
timestamp 1560284232
transform -1 0 744 0 -1 1810
box 0 0 96 200
use AOI21X1  AOI21X1_10
timestamp 1560284232
transform 1 0 744 0 -1 1810
box 0 0 64 200
use OAI21X1  OAI21X1_11
timestamp 1560284232
transform 1 0 808 0 -1 1810
box 0 0 64 200
use DFFSR  DFFSR_25
timestamp 1560284232
transform -1 0 1224 0 -1 1810
box 0 0 352 200
use BUFX2  BUFX2_5
timestamp 1560284232
transform -1 0 1272 0 -1 1810
box 0 0 48 200
use MUX2X1  MUX2X1_2
timestamp 1560284232
transform 1 0 1272 0 -1 1810
box 0 0 96 200
use INVX1  INVX1_39
timestamp 1560284232
transform -1 0 1400 0 -1 1810
box 0 0 32 200
use INVX1  INVX1_9
timestamp 1560284232
transform -1 0 1432 0 -1 1810
box 0 0 32 200
use NOR2X1  NOR2X1_3
timestamp 1560284232
transform 1 0 1432 0 -1 1810
box 0 0 48 200
use INVX1  INVX1_4
timestamp 1560284232
transform -1 0 1512 0 -1 1810
box 0 0 32 200
use FILL  FILL_8_1_0
timestamp 1560284232
transform -1 0 1528 0 -1 1810
box 0 0 16 200
use FILL  FILL_8_1_1
timestamp 1560284232
transform -1 0 1544 0 -1 1810
box 0 0 16 200
use FILL  FILL_8_1_2
timestamp 1560284232
transform -1 0 1560 0 -1 1810
box 0 0 16 200
use DFFSR  DFFSR_7
timestamp 1560284232
transform -1 0 1912 0 -1 1810
box 0 0 352 200
use DFFSR  DFFSR_24
timestamp 1560284232
transform 1 0 1912 0 -1 1810
box 0 0 352 200
use BUFX2  BUFX2_24
timestamp 1560284232
transform -1 0 56 0 1 1410
box 0 0 48 200
use DFFSR  DFFSR_29
timestamp 1560284232
transform -1 0 408 0 1 1410
box 0 0 352 200
use OAI21X1  OAI21X1_5
timestamp 1560284232
transform -1 0 472 0 1 1410
box 0 0 64 200
use AOI21X1  AOI21X1_4
timestamp 1560284232
transform -1 0 536 0 1 1410
box 0 0 64 200
use INVX1  INVX1_10
timestamp 1560284232
transform 1 0 536 0 1 1410
box 0 0 32 200
use FILL  FILL_7_0_0
timestamp 1560284232
transform 1 0 568 0 1 1410
box 0 0 16 200
use FILL  FILL_7_0_1
timestamp 1560284232
transform 1 0 584 0 1 1410
box 0 0 16 200
use FILL  FILL_7_0_2
timestamp 1560284232
transform 1 0 600 0 1 1410
box 0 0 16 200
use DFFSR  DFFSR_28
timestamp 1560284232
transform 1 0 616 0 1 1410
box 0 0 352 200
use DFFSR  DFFSR_2
timestamp 1560284232
transform 1 0 968 0 1 1410
box 0 0 352 200
use OAI21X1  OAI21X1_2
timestamp 1560284232
transform -1 0 1384 0 1 1410
box 0 0 64 200
use INVX1  INVX1_2
timestamp 1560284232
transform -1 0 1416 0 1 1410
box 0 0 32 200
use INVX1  INVX1_3
timestamp 1560284232
transform -1 0 1448 0 1 1410
box 0 0 32 200
use AND2X2  AND2X2_4
timestamp 1560284232
transform 1 0 1448 0 1 1410
box 0 0 64 200
use BUFX2  BUFX2_8
timestamp 1560284232
transform 1 0 1512 0 1 1410
box 0 0 48 200
use FILL  FILL_7_1_0
timestamp 1560284232
transform 1 0 1560 0 1 1410
box 0 0 16 200
use FILL  FILL_7_1_1
timestamp 1560284232
transform 1 0 1576 0 1 1410
box 0 0 16 200
use FILL  FILL_7_1_2
timestamp 1560284232
transform 1 0 1592 0 1 1410
box 0 0 16 200
use CLKBUF1  CLKBUF1_4
timestamp 1560284232
transform 1 0 1608 0 1 1410
box 0 0 144 200
use AOI21X1  AOI21X1_11
timestamp 1560284232
transform 1 0 1752 0 1 1410
box 0 0 64 200
use INVX1  INVX1_22
timestamp 1560284232
transform -1 0 1848 0 1 1410
box 0 0 32 200
use DFFSR  DFFSR_33
timestamp 1560284232
transform 1 0 1848 0 1 1410
box 0 0 352 200
use BUFX2  BUFX2_18
timestamp 1560284232
transform 1 0 2200 0 1 1410
box 0 0 48 200
use FILL  FILL_8_1
timestamp 1560284232
transform 1 0 2248 0 1 1410
box 0 0 16 200
use BUFX2  BUFX2_30
timestamp 1560284232
transform -1 0 56 0 -1 1410
box 0 0 48 200
use INVX1  INVX1_13
timestamp 1560284232
transform 1 0 56 0 -1 1410
box 0 0 32 200
use MUX2X1  MUX2X1_4
timestamp 1560284232
transform -1 0 184 0 -1 1410
box 0 0 96 200
use DFFSR  DFFSR_18
timestamp 1560284232
transform -1 0 536 0 -1 1410
box 0 0 352 200
use OAI21X1  OAI21X1_6
timestamp 1560284232
transform 1 0 536 0 -1 1410
box 0 0 64 200
use BUFX2  BUFX2_2
timestamp 1560284232
transform -1 0 648 0 -1 1410
box 0 0 48 200
use FILL  FILL_6_0_0
timestamp 1560284232
transform 1 0 648 0 -1 1410
box 0 0 16 200
use FILL  FILL_6_0_1
timestamp 1560284232
transform 1 0 664 0 -1 1410
box 0 0 16 200
use FILL  FILL_6_0_2
timestamp 1560284232
transform 1 0 680 0 -1 1410
box 0 0 16 200
use BUFX2  BUFX2_1
timestamp 1560284232
transform 1 0 696 0 -1 1410
box 0 0 48 200
use AOI21X1  AOI21X1_5
timestamp 1560284232
transform -1 0 808 0 -1 1410
box 0 0 64 200
use MUX2X1  MUX2X1_3
timestamp 1560284232
transform 1 0 808 0 -1 1410
box 0 0 96 200
use INVX1  INVX1_11
timestamp 1560284232
transform -1 0 936 0 -1 1410
box 0 0 32 200
use CLKBUF1  CLKBUF1_5
timestamp 1560284232
transform -1 0 1080 0 -1 1410
box 0 0 144 200
use DFFSR  DFFSR_5
timestamp 1560284232
transform 1 0 1080 0 -1 1410
box 0 0 352 200
use INVX1  INVX1_23
timestamp 1560284232
transform 1 0 1432 0 -1 1410
box 0 0 32 200
use FILL  FILL_6_1_0
timestamp 1560284232
transform 1 0 1464 0 -1 1410
box 0 0 16 200
use FILL  FILL_6_1_1
timestamp 1560284232
transform 1 0 1480 0 -1 1410
box 0 0 16 200
use FILL  FILL_6_1_2
timestamp 1560284232
transform 1 0 1496 0 -1 1410
box 0 0 16 200
use DFFSR  DFFSR_1
timestamp 1560284232
transform 1 0 1512 0 -1 1410
box 0 0 352 200
use DFFSR  DFFSR_12
timestamp 1560284232
transform 1 0 1864 0 -1 1410
box 0 0 352 200
use FILL  FILL_7_1
timestamp 1560284232
transform -1 0 2232 0 -1 1410
box 0 0 16 200
use FILL  FILL_7_2
timestamp 1560284232
transform -1 0 2248 0 -1 1410
box 0 0 16 200
use FILL  FILL_7_3
timestamp 1560284232
transform -1 0 2264 0 -1 1410
box 0 0 16 200
use BUFX2  BUFX2_33
timestamp 1560284232
transform -1 0 56 0 1 1010
box 0 0 48 200
use BUFX2  BUFX2_32
timestamp 1560284232
transform -1 0 104 0 1 1010
box 0 0 48 200
use INVX1  INVX1_14
timestamp 1560284232
transform 1 0 104 0 1 1010
box 0 0 32 200
use INVX1  INVX1_16
timestamp 1560284232
transform 1 0 136 0 1 1010
box 0 0 32 200
use AOI21X1  AOI21X1_7
timestamp 1560284232
transform 1 0 168 0 1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_8
timestamp 1560284232
transform 1 0 232 0 1 1010
box 0 0 64 200
use AOI21X1  AOI21X1_6
timestamp 1560284232
transform 1 0 296 0 1 1010
box 0 0 64 200
use DFFSR  DFFSR_20
timestamp 1560284232
transform -1 0 712 0 1 1010
box 0 0 352 200
use FILL  FILL_5_0_0
timestamp 1560284232
transform 1 0 712 0 1 1010
box 0 0 16 200
use FILL  FILL_5_0_1
timestamp 1560284232
transform 1 0 728 0 1 1010
box 0 0 16 200
use FILL  FILL_5_0_2
timestamp 1560284232
transform 1 0 744 0 1 1010
box 0 0 16 200
use INVX1  INVX1_12
timestamp 1560284232
transform 1 0 760 0 1 1010
box 0 0 32 200
use CLKBUF1  CLKBUF1_1
timestamp 1560284232
transform -1 0 936 0 1 1010
box 0 0 144 200
use DFFSR  DFFSR_3
timestamp 1560284232
transform 1 0 936 0 1 1010
box 0 0 352 200
use NAND3X1  NAND3X1_2
timestamp 1560284232
transform 1 0 1288 0 1 1010
box 0 0 64 200
use INVX1  INVX1_30
timestamp 1560284232
transform 1 0 1352 0 1 1010
box 0 0 32 200
use NOR2X1  NOR2X1_11
timestamp 1560284232
transform 1 0 1384 0 1 1010
box 0 0 48 200
use INVX1  INVX1_31
timestamp 1560284232
transform -1 0 1464 0 1 1010
box 0 0 32 200
use OAI21X1  OAI21X1_22
timestamp 1560284232
transform -1 0 1528 0 1 1010
box 0 0 64 200
use NOR2X1  NOR2X1_12
timestamp 1560284232
transform 1 0 1528 0 1 1010
box 0 0 48 200
use FILL  FILL_5_1_0
timestamp 1560284232
transform 1 0 1576 0 1 1010
box 0 0 16 200
use FILL  FILL_5_1_1
timestamp 1560284232
transform 1 0 1592 0 1 1010
box 0 0 16 200
use FILL  FILL_5_1_2
timestamp 1560284232
transform 1 0 1608 0 1 1010
box 0 0 16 200
use AOI21X1  AOI21X1_14
timestamp 1560284232
transform 1 0 1624 0 1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_25
timestamp 1560284232
transform 1 0 1688 0 1 1010
box 0 0 64 200
use AOI22X1  AOI22X1_1
timestamp 1560284232
transform -1 0 1832 0 1 1010
box 0 0 80 200
use INVX1  INVX1_1
timestamp 1560284232
transform -1 0 1864 0 1 1010
box 0 0 32 200
use BUFX2  BUFX2_15
timestamp 1560284232
transform 1 0 1864 0 1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_23
timestamp 1560284232
transform -1 0 1976 0 1 1010
box 0 0 64 200
use OAI21X1  OAI21X1_21
timestamp 1560284232
transform -1 0 2040 0 1 1010
box 0 0 64 200
use NAND2X1  NAND2X1_5
timestamp 1560284232
transform 1 0 2040 0 1 1010
box 0 0 48 200
use AOI21X1  AOI21X1_13
timestamp 1560284232
transform 1 0 2088 0 1 1010
box 0 0 64 200
use INVX1  INVX1_28
timestamp 1560284232
transform -1 0 2184 0 1 1010
box 0 0 32 200
use BUFX2  BUFX2_14
timestamp 1560284232
transform 1 0 2184 0 1 1010
box 0 0 48 200
use FILL  FILL_6_1
timestamp 1560284232
transform 1 0 2232 0 1 1010
box 0 0 16 200
use FILL  FILL_6_2
timestamp 1560284232
transform 1 0 2248 0 1 1010
box 0 0 16 200
use DFFSR  DFFSR_21
timestamp 1560284232
transform -1 0 360 0 -1 1010
box 0 0 352 200
use BUFX2  BUFX2_31
timestamp 1560284232
transform -1 0 408 0 -1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_7
timestamp 1560284232
transform -1 0 472 0 -1 1010
box 0 0 64 200
use XNOR2X1  XNOR2X1_2
timestamp 1560284232
transform -1 0 584 0 -1 1010
box 0 0 112 200
use BUFX2  BUFX2_4
timestamp 1560284232
transform -1 0 632 0 -1 1010
box 0 0 48 200
use FILL  FILL_4_0_0
timestamp 1560284232
transform -1 0 648 0 -1 1010
box 0 0 16 200
use FILL  FILL_4_0_1
timestamp 1560284232
transform -1 0 664 0 -1 1010
box 0 0 16 200
use FILL  FILL_4_0_2
timestamp 1560284232
transform -1 0 680 0 -1 1010
box 0 0 16 200
use DFFSR  DFFSR_19
timestamp 1560284232
transform -1 0 1032 0 -1 1010
box 0 0 352 200
use BUFX2  BUFX2_6
timestamp 1560284232
transform -1 0 1080 0 -1 1010
box 0 0 48 200
use BUFX2  BUFX2_9
timestamp 1560284232
transform -1 0 1128 0 -1 1010
box 0 0 48 200
use BUFX2  BUFX2_7
timestamp 1560284232
transform 1 0 1128 0 -1 1010
box 0 0 48 200
use NAND3X1  NAND3X1_7
timestamp 1560284232
transform -1 0 1240 0 -1 1010
box 0 0 64 200
use NAND3X1  NAND3X1_8
timestamp 1560284232
transform 1 0 1240 0 -1 1010
box 0 0 64 200
use INVX1  INVX1_29
timestamp 1560284232
transform -1 0 1336 0 -1 1010
box 0 0 32 200
use DFFSR  DFFSR_13
timestamp 1560284232
transform -1 0 1688 0 -1 1010
box 0 0 352 200
use FILL  FILL_4_1_0
timestamp 1560284232
transform 1 0 1688 0 -1 1010
box 0 0 16 200
use FILL  FILL_4_1_1
timestamp 1560284232
transform 1 0 1704 0 -1 1010
box 0 0 16 200
use FILL  FILL_4_1_2
timestamp 1560284232
transform 1 0 1720 0 -1 1010
box 0 0 16 200
use DFFSR  DFFSR_10
timestamp 1560284232
transform 1 0 1736 0 -1 1010
box 0 0 352 200
use NAND2X1  NAND2X1_6
timestamp 1560284232
transform -1 0 2136 0 -1 1010
box 0 0 48 200
use OAI21X1  OAI21X1_24
timestamp 1560284232
transform 1 0 2136 0 -1 1010
box 0 0 64 200
use NAND3X1  NAND3X1_6
timestamp 1560284232
transform 1 0 2200 0 -1 1010
box 0 0 64 200
use DFFSR  DFFSR_22
timestamp 1560284232
transform -1 0 360 0 1 610
box 0 0 352 200
use OAI21X1  OAI21X1_10
timestamp 1560284232
transform 1 0 360 0 1 610
box 0 0 64 200
use OAI21X1  OAI21X1_9
timestamp 1560284232
transform -1 0 488 0 1 610
box 0 0 64 200
use AOI21X1  AOI21X1_3
timestamp 1560284232
transform 1 0 488 0 1 610
box 0 0 64 200
use OAI21X1  OAI21X1_3
timestamp 1560284232
transform 1 0 552 0 1 610
box 0 0 64 200
use FILL  FILL_3_0_0
timestamp 1560284232
transform 1 0 616 0 1 610
box 0 0 16 200
use FILL  FILL_3_0_1
timestamp 1560284232
transform 1 0 632 0 1 610
box 0 0 16 200
use FILL  FILL_3_0_2
timestamp 1560284232
transform 1 0 648 0 1 610
box 0 0 16 200
use INVX1  INVX1_6
timestamp 1560284232
transform 1 0 664 0 1 610
box 0 0 32 200
use NOR2X1  NOR2X1_6
timestamp 1560284232
transform -1 0 744 0 1 610
box 0 0 48 200
use OAI21X1  OAI21X1_4
timestamp 1560284232
transform -1 0 808 0 1 610
box 0 0 64 200
use DFFSR  DFFSR_16
timestamp 1560284232
transform 1 0 808 0 1 610
box 0 0 352 200
use INVX1  INVX1_38
timestamp 1560284232
transform 1 0 1160 0 1 610
box 0 0 32 200
use INVX1  INVX1_35
timestamp 1560284232
transform -1 0 1224 0 1 610
box 0 0 32 200
use AOI22X1  AOI22X1_2
timestamp 1560284232
transform 1 0 1224 0 1 610
box 0 0 80 200
use NOR3X1  NOR3X1_1
timestamp 1560284232
transform 1 0 1304 0 1 610
box 0 0 128 200
use FILL  FILL_3_1_0
timestamp 1560284232
transform 1 0 1432 0 1 610
box 0 0 16 200
use FILL  FILL_3_1_1
timestamp 1560284232
transform 1 0 1448 0 1 610
box 0 0 16 200
use FILL  FILL_3_1_2
timestamp 1560284232
transform 1 0 1464 0 1 610
box 0 0 16 200
use DFFSR  DFFSR_11
timestamp 1560284232
transform 1 0 1480 0 1 610
box 0 0 352 200
use OAI21X1  OAI21X1_20
timestamp 1560284232
transform 1 0 1832 0 1 610
box 0 0 64 200
use OAI21X1  OAI21X1_17
timestamp 1560284232
transform 1 0 1896 0 1 610
box 0 0 64 200
use AOI21X1  AOI21X1_12
timestamp 1560284232
transform -1 0 2024 0 1 610
box 0 0 64 200
use OAI21X1  OAI21X1_16
timestamp 1560284232
transform -1 0 2088 0 1 610
box 0 0 64 200
use NAND3X1  NAND3X1_4
timestamp 1560284232
transform 1 0 2088 0 1 610
box 0 0 64 200
use OAI21X1  OAI21X1_18
timestamp 1560284232
transform 1 0 2152 0 1 610
box 0 0 64 200
use NOR2X1  NOR2X1_10
timestamp 1560284232
transform -1 0 2264 0 1 610
box 0 0 48 200
use BUFX2  BUFX2_34
timestamp 1560284232
transform -1 0 56 0 -1 610
box 0 0 48 200
use BUFX2  BUFX2_35
timestamp 1560284232
transform -1 0 104 0 -1 610
box 0 0 48 200
use MUX2X1  MUX2X1_6
timestamp 1560284232
transform -1 0 200 0 -1 610
box 0 0 96 200
use INVX1  INVX1_18
timestamp 1560284232
transform -1 0 232 0 -1 610
box 0 0 32 200
use AOI21X1  AOI21X1_8
timestamp 1560284232
transform 1 0 232 0 -1 610
box 0 0 64 200
use AOI21X1  AOI21X1_9
timestamp 1560284232
transform 1 0 296 0 -1 610
box 0 0 64 200
use INVX1  INVX1_20
timestamp 1560284232
transform -1 0 392 0 -1 610
box 0 0 32 200
use XNOR2X1  XNOR2X1_1
timestamp 1560284232
transform -1 0 504 0 -1 610
box 0 0 112 200
use MUX2X1  MUX2X1_7
timestamp 1560284232
transform 1 0 504 0 -1 610
box 0 0 96 200
use BUFX2  BUFX2_3
timestamp 1560284232
transform -1 0 648 0 -1 610
box 0 0 48 200
use FILL  FILL_2_0_0
timestamp 1560284232
transform -1 0 664 0 -1 610
box 0 0 16 200
use FILL  FILL_2_0_1
timestamp 1560284232
transform -1 0 680 0 -1 610
box 0 0 16 200
use FILL  FILL_2_0_2
timestamp 1560284232
transform -1 0 696 0 -1 610
box 0 0 16 200
use INVX1  INVX1_19
timestamp 1560284232
transform -1 0 728 0 -1 610
box 0 0 32 200
use CLKBUF1  CLKBUF1_2
timestamp 1560284232
transform -1 0 872 0 -1 610
box 0 0 144 200
use CLKBUF1  CLKBUF1_3
timestamp 1560284232
transform 1 0 872 0 -1 610
box 0 0 144 200
use NOR2X1  NOR2X1_14
timestamp 1560284232
transform 1 0 1016 0 -1 610
box 0 0 48 200
use NAND2X1  NAND2X1_7
timestamp 1560284232
transform -1 0 1112 0 -1 610
box 0 0 48 200
use NAND3X1  NAND3X1_1
timestamp 1560284232
transform 1 0 1112 0 -1 610
box 0 0 64 200
use NAND3X1  NAND3X1_5
timestamp 1560284232
transform -1 0 1240 0 -1 610
box 0 0 64 200
use DFFSR  DFFSR_14
timestamp 1560284232
transform -1 0 1592 0 -1 610
box 0 0 352 200
use FILL  FILL_2_1_0
timestamp 1560284232
transform 1 0 1592 0 -1 610
box 0 0 16 200
use FILL  FILL_2_1_1
timestamp 1560284232
transform 1 0 1608 0 -1 610
box 0 0 16 200
use FILL  FILL_2_1_2
timestamp 1560284232
transform 1 0 1624 0 -1 610
box 0 0 16 200
use OAI21X1  OAI21X1_28
timestamp 1560284232
transform 1 0 1640 0 -1 610
box 0 0 64 200
use AND2X2  AND2X2_2
timestamp 1560284232
transform 1 0 1704 0 -1 610
box 0 0 64 200
use OAI21X1  OAI21X1_19
timestamp 1560284232
transform -1 0 1832 0 -1 610
box 0 0 64 200
use NOR2X1  NOR2X1_1
timestamp 1560284232
transform -1 0 1880 0 -1 610
box 0 0 48 200
use XOR2X1  XOR2X1_1
timestamp 1560284232
transform 1 0 1880 0 -1 610
box 0 0 112 200
use OAI21X1  OAI21X1_14
timestamp 1560284232
transform -1 0 2056 0 -1 610
box 0 0 64 200
use BUFX2  BUFX2_12
timestamp 1560284232
transform 1 0 2056 0 -1 610
box 0 0 48 200
use INVX1  INVX1_25
timestamp 1560284232
transform 1 0 2104 0 -1 610
box 0 0 32 200
use NOR2X1  NOR2X1_8
timestamp 1560284232
transform 1 0 2136 0 -1 610
box 0 0 48 200
use NAND2X1  NAND2X1_2
timestamp 1560284232
transform -1 0 2232 0 -1 610
box 0 0 48 200
use FILL  FILL_3_1
timestamp 1560284232
transform -1 0 2248 0 -1 610
box 0 0 16 200
use FILL  FILL_3_2
timestamp 1560284232
transform -1 0 2264 0 -1 610
box 0 0 16 200
use INVX1  INVX1_17
timestamp 1560284232
transform 1 0 8 0 1 210
box 0 0 32 200
use DFFSR  DFFSR_23
timestamp 1560284232
transform -1 0 392 0 1 210
box 0 0 352 200
use DFFSR  DFFSR_4
timestamp 1560284232
transform 1 0 392 0 1 210
box 0 0 352 200
use FILL  FILL_1_0_0
timestamp 1560284232
transform 1 0 744 0 1 210
box 0 0 16 200
use FILL  FILL_1_0_1
timestamp 1560284232
transform 1 0 760 0 1 210
box 0 0 16 200
use FILL  FILL_1_0_2
timestamp 1560284232
transform 1 0 776 0 1 210
box 0 0 16 200
use NAND2X1  NAND2X1_1
timestamp 1560284232
transform 1 0 792 0 1 210
box 0 0 48 200
use OAI21X1  OAI21X1_1
timestamp 1560284232
transform -1 0 904 0 1 210
box 0 0 64 200
use OAI21X1  OAI21X1_30
timestamp 1560284232
transform 1 0 904 0 1 210
box 0 0 64 200
use INVX1  INVX1_37
timestamp 1560284232
transform 1 0 968 0 1 210
box 0 0 32 200
use NAND3X1  NAND3X1_11
timestamp 1560284232
transform 1 0 1000 0 1 210
box 0 0 64 200
use NAND3X1  NAND3X1_12
timestamp 1560284232
transform -1 0 1128 0 1 210
box 0 0 64 200
use AND2X2  AND2X2_3
timestamp 1560284232
transform -1 0 1192 0 1 210
box 0 0 64 200
use NOR2X1  NOR2X1_2
timestamp 1560284232
transform 1 0 1192 0 1 210
box 0 0 48 200
use DFFSR  DFFSR_8
timestamp 1560284232
transform -1 0 1592 0 1 210
box 0 0 352 200
use FILL  FILL_1_1_0
timestamp 1560284232
transform 1 0 1592 0 1 210
box 0 0 16 200
use FILL  FILL_1_1_1
timestamp 1560284232
transform 1 0 1608 0 1 210
box 0 0 16 200
use FILL  FILL_1_1_2
timestamp 1560284232
transform 1 0 1624 0 1 210
box 0 0 16 200
use INVX1  INVX1_26
timestamp 1560284232
transform 1 0 1640 0 1 210
box 0 0 32 200
use NAND2X1  NAND2X1_3
timestamp 1560284232
transform 1 0 1672 0 1 210
box 0 0 48 200
use NOR2X1  NOR2X1_9
timestamp 1560284232
transform -1 0 1768 0 1 210
box 0 0 48 200
use INVX1  INVX1_27
timestamp 1560284232
transform 1 0 1768 0 1 210
box 0 0 32 200
use OAI21X1  OAI21X1_15
timestamp 1560284232
transform 1 0 1800 0 1 210
box 0 0 64 200
use NAND2X1  NAND2X1_4
timestamp 1560284232
transform -1 0 1912 0 1 210
box 0 0 48 200
use NAND3X1  NAND3X1_10
timestamp 1560284232
transform 1 0 1912 0 1 210
box 0 0 64 200
use OAI21X1  OAI21X1_26
timestamp 1560284232
transform -1 0 2040 0 1 210
box 0 0 64 200
use INVX1  INVX1_34
timestamp 1560284232
transform 1 0 2040 0 1 210
box 0 0 32 200
use OAI21X1  OAI21X1_27
timestamp 1560284232
transform -1 0 2136 0 1 210
box 0 0 64 200
use NAND3X1  NAND3X1_9
timestamp 1560284232
transform 1 0 2136 0 1 210
box 0 0 64 200
use NOR2X1  NOR2X1_13
timestamp 1560284232
transform 1 0 2200 0 1 210
box 0 0 48 200
use FILL  FILL_2_1
timestamp 1560284232
transform 1 0 2248 0 1 210
box 0 0 16 200
use BUFX2  BUFX2_26
timestamp 1560284232
transform -1 0 56 0 -1 210
box 0 0 48 200
use DFFSR  DFFSR_31
timestamp 1560284232
transform -1 0 408 0 -1 210
box 0 0 352 200
use DFFSR  DFFSR_32
timestamp 1560284232
transform 1 0 408 0 -1 210
box 0 0 352 200
use FILL  FILL_0_0_0
timestamp 1560284232
transform 1 0 760 0 -1 210
box 0 0 16 200
use FILL  FILL_0_0_1
timestamp 1560284232
transform 1 0 776 0 -1 210
box 0 0 16 200
use FILL  FILL_0_0_2
timestamp 1560284232
transform 1 0 792 0 -1 210
box 0 0 16 200
use BUFX2  BUFX2_27
timestamp 1560284232
transform 1 0 808 0 -1 210
box 0 0 48 200
use BUFX2  BUFX2_17
timestamp 1560284232
transform -1 0 904 0 -1 210
box 0 0 48 200
use DFFSR  DFFSR_15
timestamp 1560284232
transform -1 0 1256 0 -1 210
box 0 0 352 200
use BUFX2  BUFX2_16
timestamp 1560284232
transform 1 0 1256 0 -1 210
box 0 0 48 200
use BUFX2  BUFX2_10
timestamp 1560284232
transform 1 0 1304 0 -1 210
box 0 0 48 200
use NOR2X1  NOR2X1_7
timestamp 1560284232
transform 1 0 1352 0 -1 210
box 0 0 48 200
use AND2X2  AND2X2_1
timestamp 1560284232
transform 1 0 1400 0 -1 210
box 0 0 64 200
use OAI21X1  OAI21X1_12
timestamp 1560284232
transform 1 0 1464 0 -1 210
box 0 0 64 200
use OAI21X1  OAI21X1_13
timestamp 1560284232
transform -1 0 1592 0 -1 210
box 0 0 64 200
use FILL  FILL_0_1_0
timestamp 1560284232
transform -1 0 1608 0 -1 210
box 0 0 16 200
use FILL  FILL_0_1_1
timestamp 1560284232
transform -1 0 1624 0 -1 210
box 0 0 16 200
use FILL  FILL_0_1_2
timestamp 1560284232
transform -1 0 1640 0 -1 210
box 0 0 16 200
use BUFX2  BUFX2_11
timestamp 1560284232
transform -1 0 1688 0 -1 210
box 0 0 48 200
use DFFSR  DFFSR_9
timestamp 1560284232
transform -1 0 2040 0 -1 210
box 0 0 352 200
use OAI21X1  OAI21X1_29
timestamp 1560284232
transform 1 0 2040 0 -1 210
box 0 0 64 200
use INVX1  INVX1_24
timestamp 1560284232
transform -1 0 2136 0 -1 210
box 0 0 32 200
use INVX1  INVX1_36
timestamp 1560284232
transform -1 0 2168 0 -1 210
box 0 0 32 200
use INVX1  INVX1_33
timestamp 1560284232
transform -1 0 2200 0 -1 210
box 0 0 32 200
use BUFX2  BUFX2_13
timestamp 1560284232
transform 1 0 2200 0 -1 210
box 0 0 48 200
use FILL  FILL_1_1
timestamp 1560284232
transform -1 0 2264 0 -1 210
box 0 0 16 200
<< labels >>
flabel metal4 s 632 -40 680 -16 7 FreeSans 24 270 0 0 vdd
port 0 nsew
flabel metal4 s 1544 -40 1592 -16 7 FreeSans 24 270 0 0 gnd
port 1 nsew
flabel metal2 s 1629 2037 1635 2043 3 FreeSans 24 90 0 0 clock
port 2 nsew
flabel metal2 s 1373 2037 1379 2043 3 FreeSans 24 90 0 0 reset
port 3 nsew
flabel metal2 s 1821 2037 1827 2043 3 FreeSans 24 90 0 0 start
port 4 nsew
flabel metal2 s 2029 2037 2035 2043 3 FreeSans 24 90 0 0 N[0]
port 5 nsew
flabel metal3 s 2285 577 2291 583 3 FreeSans 24 0 0 0 N[1]
port 6 nsew
flabel metal3 s 2285 537 2291 543 3 FreeSans 24 0 0 0 N[2]
port 7 nsew
flabel metal3 s 2285 677 2291 683 3 FreeSans 24 0 0 0 N[3]
port 8 nsew
flabel metal3 s 2285 717 2291 723 3 FreeSans 24 0 0 0 N[4]
port 9 nsew
flabel metal3 s 2285 257 2291 263 3 FreeSans 24 0 0 0 N[5]
port 10 nsew
flabel metal3 s 2285 337 2291 343 3 FreeSans 24 0 0 0 N[6]
port 11 nsew
flabel metal3 s 2285 1857 2291 1863 3 FreeSans 24 0 0 0 N[7]
port 12 nsew
flabel metal3 s 2285 297 2291 303 3 FreeSans 24 0 0 0 N[8]
port 13 nsew
flabel metal2 s 2173 2037 2179 2043 3 FreeSans 24 90 0 0 dp[0]
port 14 nsew
flabel metal2 s 861 2037 867 2043 3 FreeSans 24 90 0 0 dp[1]
port 15 nsew
flabel metal2 s 429 2037 435 2043 3 FreeSans 24 90 0 0 dp[2]
port 16 nsew
flabel metal2 s 1597 2037 1603 2043 3 FreeSans 24 90 0 0 dp[3]
port 17 nsew
flabel metal2 s 973 2037 979 2043 3 FreeSans 24 90 0 0 dp[4]
port 18 nsew
flabel metal3 s -19 1497 -13 1503 7 FreeSans 24 0 0 0 dp[5]
port 19 nsew
flabel metal3 s -19 1897 -13 1903 7 FreeSans 24 0 0 0 dp[6]
port 20 nsew
flabel metal3 s -19 97 -13 103 7 FreeSans 24 0 0 0 dp[7]
port 21 nsew
flabel metal2 s 813 -23 819 -17 7 FreeSans 24 270 0 0 dp[8]
port 22 nsew
flabel metal3 s 2285 1497 2291 1503 3 FreeSans 24 0 0 0 done
port 23 nsew
flabel metal2 s 1325 -23 1331 -17 7 FreeSans 24 270 0 0 counter[0]
port 24 nsew
flabel metal2 s 1661 -23 1667 -17 7 FreeSans 24 270 0 0 counter[1]
port 25 nsew
flabel metal3 s 2285 497 2291 503 3 FreeSans 24 0 0 0 counter[2]
port 26 nsew
flabel metal3 s 2285 97 2291 103 3 FreeSans 24 0 0 0 counter[3]
port 27 nsew
flabel metal3 s 2285 1137 2291 1143 3 FreeSans 24 0 0 0 counter[4]
port 28 nsew
flabel metal3 s 2285 1097 2291 1103 3 FreeSans 24 0 0 0 counter[5]
port 29 nsew
flabel metal2 s 1277 -23 1283 -17 7 FreeSans 24 270 0 0 counter[6]
port 30 nsew
flabel metal2 s 877 -23 883 -17 7 FreeSans 24 270 0 0 counter[7]
port 31 nsew
flabel metal2 s 925 2037 931 2043 3 FreeSans 24 90 0 0 sr[0]
port 32 nsew
flabel metal3 s -19 1697 -13 1703 7 FreeSans 24 0 0 0 sr[1]
port 33 nsew
flabel metal3 s -19 1297 -13 1303 7 FreeSans 24 0 0 0 sr[2]
port 34 nsew
flabel metal3 s -19 897 -13 903 7 FreeSans 24 0 0 0 sr[3]
port 35 nsew
flabel metal3 s -19 1097 -13 1103 7 FreeSans 24 0 0 0 sr[4]
port 36 nsew
flabel metal3 s -19 1137 -13 1143 7 FreeSans 24 0 0 0 sr[5]
port 37 nsew
flabel metal3 s -19 537 -13 543 7 FreeSans 24 0 0 0 sr[6]
port 38 nsew
flabel metal3 s -19 497 -13 503 7 FreeSans 24 0 0 0 sr[7]
port 39 nsew
<< end >>
