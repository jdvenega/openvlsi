magic
tech scmos
magscale 1 2
timestamp 1556508158
<< checkpaint >>
rect -78 -66 134 270
<< nwell >>
rect -18 96 74 210
<< ntransistor >>
rect 14 12 18 42
rect 30 12 34 52
rect 46 12 50 52
<< ptransistor >>
rect 14 128 18 188
rect 30 108 34 188
rect 46 108 50 188
<< ndiffusion >>
rect 20 51 30 52
rect 4 41 14 42
rect 12 13 14 41
rect 4 12 14 13
rect 18 13 20 42
rect 28 13 30 51
rect 18 12 30 13
rect 34 51 46 52
rect 34 13 36 51
rect 44 13 46 51
rect 34 12 46 13
rect 50 51 60 52
rect 50 13 52 51
rect 50 12 60 13
<< pdiffusion >>
rect 4 187 14 188
rect 12 129 14 187
rect 4 128 14 129
rect 18 128 20 188
rect 28 120 30 188
rect 20 108 30 120
rect 34 187 46 188
rect 34 109 36 187
rect 44 109 46 187
rect 34 108 46 109
rect 50 187 60 188
rect 50 109 52 187
rect 50 108 60 109
<< ndcontact >>
rect 4 13 12 41
rect 20 13 28 51
rect 36 13 44 51
rect 52 13 60 51
<< pdcontact >>
rect 4 129 12 187
rect 20 120 28 188
rect 36 109 44 187
rect 52 109 60 187
<< psubstratepcontact >>
rect -4 -4 4 4
rect 28 -4 36 4
<< nsubstratencontact >>
rect -4 196 4 204
rect 28 196 36 204
<< polysilicon >>
rect 14 188 18 192
rect 30 188 34 192
rect 46 188 50 192
rect 14 42 18 128
rect 30 106 34 108
rect 46 106 50 108
rect 30 102 50 106
rect 30 88 34 102
rect 30 58 34 80
rect 30 54 50 58
rect 30 52 34 54
rect 46 52 50 54
rect 14 8 18 12
rect 30 8 34 12
rect 46 8 50 12
<< polycontact >>
rect 6 78 14 86
rect 26 80 34 88
<< metal1 >>
rect -4 204 68 206
rect 4 196 28 204
rect 36 196 68 204
rect -4 194 68 196
rect 20 188 28 194
rect 4 187 12 188
rect 4 114 12 129
rect 36 187 44 188
rect 4 108 30 114
rect 52 187 60 194
rect 44 109 46 118
rect 36 108 46 109
rect 52 108 60 109
rect 4 86 14 94
rect 24 88 30 108
rect 24 80 26 88
rect 24 64 30 80
rect 40 74 46 108
rect 36 66 46 74
rect 4 58 30 64
rect 4 41 12 58
rect 40 52 46 66
rect 4 12 12 13
rect 20 51 28 52
rect 20 6 28 13
rect 36 51 46 52
rect 44 46 46 51
rect 52 51 60 52
rect 36 12 44 13
rect 52 6 60 13
rect -4 4 68 6
rect 4 -4 28 4
rect 36 -4 68 4
rect -4 -6 68 -4
<< m1p >>
rect 4 86 12 94
rect 36 66 44 74
<< labels >>
rlabel metal1 8 200 8 200 4 vdd
rlabel metal1 8 0 8 0 4 gnd
rlabel metal1 8 90 8 90 4 A
rlabel metal1 40 70 40 70 4 Y
<< properties >>
string path 18.000 33.000 22.000 33.000 22.000 37.000 18.000 37.000 18.000 33.000 
<< end >>
